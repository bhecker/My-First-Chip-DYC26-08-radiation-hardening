* NGSPICE file created from top.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_IOPadIn abstract view
.subckt sg13g2_IOPadIn iovdd iovss p2c pad vdd vss
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_Filler200 abstract view
.subckt sg13g2_Filler200 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_Filler400 abstract view
.subckt sg13g2_Filler400 iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for bondpad_70x70 abstract view
.subckt bondpad_70x70 pad
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_IOPadOut30mA abstract view
.subckt sg13g2_IOPadOut30mA c2p iovdd iovss pad vdd vss
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_Corner abstract view
.subckt sg13g2_Corner iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_16 abstract view
.subckt sg13g2_buf_16 X A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_IOPadVss abstract view
.subckt sg13g2_IOPadVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVss abstract view
.subckt sg13g2_IOPadIOVss iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadIOVdd abstract view
.subckt sg13g2_IOPadIOVdd iovdd iovss vdd vss
.ends

* Black-box entry subcircuit for sg13g2_IOPadVdd abstract view
.subckt sg13g2_IOPadVdd iovdd iovss vdd vss
.ends

.subckt top IOVDD IOVSS VDD VSS clk_PAD in_data_PADs[0] in_data_PADs[1] in_data_PADs[2]
+ in_data_PADs[3] in_data_PADs[4] in_data_PADs[5] in_data_PADs[6] in_data_PADs[7]
+ in_ready_PAD in_valid_PAD out_data_PADs[0] out_data_PADs[1] out_data_PADs[2] out_data_PADs[3]
+ out_data_PADs[4] out_data_PADs[5] out_data_PADs[6] out_data_PADs[7] out_ready_PAD
+ out_valid_PAD rst_n_PAD
XFILLER_79_391 VDD VSS sg13g2_decap_8
XFILLER_67_553 VDD VSS sg13g2_decap_8
XFILLER_54_203 VDD VSS sg13g2_decap_8
XFILLER_27_406 VDD VSS sg13g2_decap_8
XFILLER_39_266 VDD VSS sg13g2_decap_8
XFILLER_82_534 VDD VSS sg13g2_decap_8
XFILLER_55_748 VDD VSS sg13g2_decap_8
XFILLER_54_214 VDD VSS sg13g2_fill_2
X_2106_ _2106_/A _2106_/B _2106_/C _2106_/Y VDD VSS sg13g2_nor3_1
X_2037_ _2037_/A _2037_/B _2037_/X VDD VSS sg13g2_and2_1
XFILLER_36_973 VDD VSS sg13g2_decap_8
XFILLER_51_932 VDD VSS sg13g2_decap_8
XFILLER_23_623 VDD VSS sg13g2_decap_8
XFILLER_35_483 VDD VSS sg13g2_decap_8
XFILLER_62_280 VDD VSS sg13g2_decap_8
XFILLER_22_133 VDD VSS sg13g2_decap_8
XFILLER_50_486 VDD VSS sg13g2_decap_4
XFILLER_50_497 VDD VSS sg13g2_decap_8
XFILLER_109_728 VDD VSS sg13g2_decap_8
XFILLER_105_945 VDD VSS sg13g2_decap_8
Xhold362 _2193_/Q VDD VSS hold362/X sg13g2_dlygate4sd3_1
Xhold351 _2177_/Q VDD VSS hold351/X sg13g2_dlygate4sd3_1
Xhold340 _2264_/Q VDD VSS _1487_/A sg13g2_dlygate4sd3_1
XFILLER_7_7 VDD VSS sg13g2_decap_8
XFILLER_81_1029 VDD VSS sg13g2_fill_1
XFILLER_104_444 VDD VSS sg13g2_decap_8
XFILLER_89_133 VDD VSS sg13g2_decap_8
Xhold395 _1268_/Y VDD VSS _1269_/A sg13g2_dlygate4sd3_1
Xhold384 _1310_/Y VDD VSS _1311_/A sg13g2_dlygate4sd3_1
Xhold373 _2255_/Q VDD VSS _1198_/A sg13g2_dlygate4sd3_1
X_2205__130 VDD VSS _2205_/RESET_B sg13g2_tiehi
XFILLER_100_661 VDD VSS sg13g2_decap_8
XFILLER_86_862 VDD VSS sg13g2_decap_8
XFILLER_93_14 VDD VSS sg13g2_decap_8
XFILLER_46_726 VDD VSS sg13g2_decap_8
XFILLER_18_406 VDD VSS sg13g2_decap_8
XFILLER_73_545 VDD VSS sg13g2_decap_8
XFILLER_85_383 VDD VSS sg13g2_decap_8
XFILLER_45_203 VDD VSS sg13g2_decap_8
XFILLER_73_556 VDD VSS sg13g2_fill_1
XFILLER_73_567 VDD VSS sg13g2_decap_8
XFILLER_27_973 VDD VSS sg13g2_decap_8
XFILLER_61_707 VDD VSS sg13g2_decap_8
XFILLER_45_269 VDD VSS sg13g2_decap_8
XFILLER_42_910 VDD VSS sg13g2_decap_8
XFILLER_60_228 VDD VSS sg13g2_decap_8
XFILLER_14_623 VDD VSS sg13g2_decap_8
XFILLER_26_63 VDD VSS sg13g2_decap_8
XFILLER_26_483 VDD VSS sg13g2_decap_8
XFILLER_13_133 VDD VSS sg13g2_decap_8
XFILLER_42_987 VDD VSS sg13g2_decap_8
XFILLER_9_126 VDD VSS sg13g2_decap_8
XFILLER_10_840 VDD VSS sg13g2_decap_8
XFILLER_42_84 VDD VSS sg13g2_decap_8
XFILLER_6_833 VDD VSS sg13g2_decap_8
XFILLER_5_343 VDD VSS sg13g2_decap_8
XFILLER_108_794 VDD VSS sg13g2_decap_8
XFILLER_96_637 VDD VSS sg13g2_decap_8
XFILLER_110_403 VDD VSS sg13g2_decap_8
XFILLER_3_56 VDD VSS sg13g2_decap_8
XFILLER_1_560 VDD VSS sg13g2_decap_8
XFILLER_111_959 VDD VSS sg13g2_decap_8
X_1270_ _1270_/Y _1280_/B1 hold325/X _1280_/A2 _2315_/Q VDD VSS sg13g2_a22oi_1
XFILLER_77_851 VDD VSS sg13g2_fill_1
XFILLER_95_147 VDD VSS sg13g2_decap_8
XFILLER_77_884 VDD VSS sg13g2_decap_8
XFILLER_76_350 VDD VSS sg13g2_decap_8
XFILLER_67_70 VDD VSS sg13g2_decap_8
XFILLER_97_1036 VDD VSS sg13g2_decap_8
XFILLER_76_394 VDD VSS sg13g2_decap_8
XFILLER_49_586 VDD VSS sg13g2_fill_2
XFILLER_3_1029 VDD VSS sg13g2_decap_8
XFILLER_36_203 VDD VSS sg13g2_decap_8
XFILLER_92_854 VDD VSS sg13g2_decap_8
XFILLER_64_578 VDD VSS sg13g2_decap_8
XFILLER_18_973 VDD VSS sg13g2_decap_8
XFILLER_91_375 VDD VSS sg13g2_decap_8
XFILLER_33_910 VDD VSS sg13g2_decap_8
XFILLER_17_483 VDD VSS sg13g2_decap_8
XFILLER_83_91 VDD VSS sg13g2_decap_8
XFILLER_32_420 VDD VSS sg13g2_decap_8
XFILLER_33_987 VDD VSS sg13g2_decap_8
XFILLER_20_637 VDD VSS sg13g2_decap_8
XFILLER_32_497 VDD VSS sg13g2_decap_8
XFILLER_9_693 VDD VSS sg13g2_decap_8
XFILLER_66_0 VDD VSS sg13g2_decap_8
XFILLER_105_208 VDD VSS sg13g2_decap_8
X_2187__166 VDD VSS _2187_/RESET_B sg13g2_tiehi
X_1606_ _1618_/A _1606_/A _1606_/B VDD VSS sg13g2_xnor2_1
XFILLER_99_442 VDD VSS sg13g2_fill_1
XFILLER_87_637 VDD VSS sg13g2_decap_8
XFILLER_99_497 VDD VSS sg13g2_decap_8
X_1537_ VSS VDD _1556_/S0 _1214_/Y _1537_/Y _1523_/B sg13g2_a21oi_1
XFILLER_59_328 VDD VSS sg13g2_fill_1
XFILLER_59_317 VDD VSS sg13g2_decap_8
X_1468_ _1367_/A VDD _1468_/Y VSS _1370_/A _1481_/A2 sg13g2_o21ai_1
X_2298__117 VDD VSS _2298_/RESET_B sg13g2_tiehi
XFILLER_110_970 VDD VSS sg13g2_decap_8
XFILLER_101_458 VDD VSS sg13g2_decap_8
X_1399_ _1400_/A _1392_/Y hold483/X _1392_/B _1376_/A VDD VSS sg13g2_a22oi_1
XFILLER_41_1035 VDD VSS sg13g2_decap_8
XFILLER_68_862 VDD VSS sg13g2_decap_8
XFILLER_67_350 VDD VSS sg13g2_decap_8
XFILLER_55_501 VDD VSS sg13g2_decap_8
X_2339__147 VDD VSS _2339_/RESET_B sg13g2_tiehi
XFILLER_67_394 VDD VSS sg13g2_decap_8
XFILLER_67_372 VDD VSS sg13g2_decap_4
XFILLER_27_203 VDD VSS sg13g2_decap_8
XFILLER_82_342 VDD VSS sg13g2_decap_8
XFILLER_103_35 VDD VSS sg13g2_decap_8
XFILLER_55_567 VDD VSS sg13g2_decap_8
XFILLER_36_770 VDD VSS sg13g2_decap_8
XFILLER_24_910 VDD VSS sg13g2_decap_8
XFILLER_63_28 VDD VSS sg13g2_decap_8
XFILLER_23_420 VDD VSS sg13g2_decap_8
XFILLER_35_280 VDD VSS sg13g2_decap_8
XFILLER_24_987 VDD VSS sg13g2_decap_8
XFILLER_51_751 VDD VSS sg13g2_decap_8
XFILLER_11_637 VDD VSS sg13g2_decap_8
XFILLER_23_497 VDD VSS sg13g2_decap_8
XFILLER_50_283 VDD VSS sg13g2_decap_8
XFILLER_10_147 VDD VSS sg13g2_decap_8
XFILLER_12_21 VDD VSS sg13g2_decap_8
XFILLER_109_525 VDD VSS sg13g2_decap_8
XFILLER_88_14 VDD VSS sg13g2_decap_8
XFILLER_12_98 VDD VSS sg13g2_decap_8
XFILLER_3_847 VDD VSS sg13g2_decap_8
XFILLER_105_742 VDD VSS sg13g2_decap_8
XFILLER_2_357 VDD VSS sg13g2_decap_8
XFILLER_104_252 VDD VSS sg13g2_decap_8
XFILLER_78_659 VDD VSS sg13g2_decap_8
XFILLER_77_147 VDD VSS sg13g2_decap_8
XFILLER_101_970 VDD VSS sg13g2_decap_8
XFILLER_93_607 VDD VSS sg13g2_decap_8
XFILLER_74_821 VDD VSS sg13g2_decap_8
XFILLER_92_117 VDD VSS sg13g2_decap_4
XFILLER_58_372 VDD VSS sg13g2_decap_4
XFILLER_18_203 VDD VSS sg13g2_decap_8
XFILLER_100_491 VDD VSS sg13g2_fill_1
XFILLER_34_707 VDD VSS sg13g2_decap_8
XFILLER_37_84 VDD VSS sg13g2_decap_8
XFILLER_74_898 VDD VSS sg13g2_decap_8
XFILLER_73_386 VDD VSS sg13g2_decap_8
XFILLER_27_770 VDD VSS sg13g2_decap_8
XFILLER_61_515 VDD VSS sg13g2_decap_8
XFILLER_15_910 VDD VSS sg13g2_decap_8
XFILLER_33_217 VDD VSS sg13g2_decap_8
X_2253__245 VDD VSS _2253_/RESET_B sg13g2_tiehi
XFILLER_57_1053 VDD VSS sg13g2_decap_8
XFILLER_57_1031 VDD VSS sg13g2_decap_4
XFILLER_14_420 VDD VSS sg13g2_decap_8
XFILLER_26_280 VDD VSS sg13g2_decap_8
XFILLER_30_924 VDD VSS sg13g2_decap_8
XFILLER_15_987 VDD VSS sg13g2_decap_8
XFILLER_18_1015 VDD VSS sg13g2_decap_8
XFILLER_42_784 VDD VSS sg13g2_decap_8
XFILLER_14_497 VDD VSS sg13g2_decap_8
XFILLER_53_83 VDD VSS sg13g2_decap_4
XFILLER_105_1029 VDD VSS sg13g2_decap_8
XFILLER_41_294 VDD VSS sg13g2_decap_8
XFILLER_6_630 VDD VSS sg13g2_decap_8
XFILLER_5_140 VDD VSS sg13g2_decap_8
XFILLER_108_591 VDD VSS sg13g2_decap_8
XFILLER_97_902 VDD VSS sg13g2_decap_8
X_2371_ _2371_/RESET_B VSS VDD _2371_/D _2371_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_64_1035 VDD VSS sg13g2_decap_8
XFILLER_68_103 VDD VSS sg13g2_decap_8
XFILLER_111_756 VDD VSS sg13g2_decap_8
X_1322_ _1322_/Y _1322_/B1 hold304/X _1322_/A2 _2324_/Q VDD VSS sg13g2_a22oi_1
XFILLER_96_434 VDD VSS sg13g2_decap_8
XFILLER_78_91 VDD VSS sg13g2_decap_8
XFILLER_25_1008 VDD VSS sg13g2_decap_8
XFILLER_110_266 VDD VSS sg13g2_decap_8
X_1253_ _1501_/A _1252_/Y _1265_/B VDD VSS sg13g2_nor2b_1
XFILLER_68_169 VDD VSS sg13g2_decap_8
XFILLER_77_681 VDD VSS sg13g2_decap_8
XFILLER_37_567 VDD VSS sg13g2_decap_8
XFILLER_25_707 VDD VSS sg13g2_decap_8
XFILLER_91_150 VDD VSS sg13g2_decap_8
XFILLER_52_526 VDD VSS sg13g2_decap_8
XFILLER_18_770 VDD VSS sg13g2_decap_8
XFILLER_24_217 VDD VSS sg13g2_decap_8
XFILLER_80_846 VDD VSS sg13g2_decap_4
XFILLER_17_280 VDD VSS sg13g2_decap_8
XFILLER_21_924 VDD VSS sg13g2_decap_8
XFILLER_33_784 VDD VSS sg13g2_decap_8
XFILLER_20_434 VDD VSS sg13g2_decap_8
XFILLER_32_294 VDD VSS sg13g2_decap_8
XFILLER_9_490 VDD VSS sg13g2_decap_8
XFILLER_106_539 VDD VSS sg13g2_decap_4
XFILLER_59_103 VDD VSS sg13g2_decap_8
XFILLER_102_756 VDD VSS sg13g2_fill_1
XFILLER_87_423 VDD VSS sg13g2_decap_8
XFILLER_88_979 VDD VSS sg13g2_decap_8
XFILLER_102_789 VDD VSS sg13g2_fill_1
XFILLER_101_255 VDD VSS sg13g2_decap_8
XFILLER_87_489 VDD VSS sg13g2_decap_4
XFILLER_83_640 VDD VSS sg13g2_decap_8
XFILLER_74_49 VDD VSS sg13g2_decap_8
XFILLER_56_843 VDD VSS sg13g2_decap_8
XFILLER_28_567 VDD VSS sg13g2_decap_8
XFILLER_16_707 VDD VSS sg13g2_decap_8
XFILLER_83_684 VDD VSS sg13g2_decap_8
XFILLER_15_217 VDD VSS sg13g2_decap_8
X_2317__242 VDD VSS _2317_/RESET_B sg13g2_tiehi
XFILLER_70_334 VDD VSS sg13g2_fill_1
XFILLER_43_559 VDD VSS sg13g2_decap_4
XFILLER_24_784 VDD VSS sg13g2_decap_8
XFILLER_12_924 VDD VSS sg13g2_decap_8
XFILLER_11_434 VDD VSS sg13g2_decap_8
XFILLER_8_917 VDD VSS sg13g2_decap_8
XFILLER_23_42 VDD VSS sg13g2_decap_8
XFILLER_23_294 VDD VSS sg13g2_decap_8
XFILLER_7_427 VDD VSS sg13g2_decap_8
XFILLER_109_333 VDD VSS sg13g2_decap_8
XFILLER_99_35 VDD VSS sg13g2_decap_8
XFILLER_109_399 VDD VSS sg13g2_decap_8
XFILLER_79_902 VDD VSS sg13g2_fill_1
XFILLER_3_644 VDD VSS sg13g2_decap_8
XFILLER_2_154 VDD VSS sg13g2_decap_8
XFILLER_79_968 VDD VSS sg13g2_decap_8
XFILLER_94_927 VDD VSS sg13g2_decap_8
XFILLER_78_478 VDD VSS sg13g2_decap_8
XFILLER_87_990 VDD VSS sg13g2_decap_8
XFILLER_78_489 VDD VSS sg13g2_fill_1
XFILLER_59_692 VDD VSS sg13g2_fill_2
XFILLER_47_810 VDD VSS sg13g2_decap_8
XFILLER_111_1022 VDD VSS sg13g2_decap_8
XFILLER_58_180 VDD VSS sg13g2_decap_8
XFILLER_0_35 VDD VSS sg13g2_decap_8
XFILLER_73_150 VDD VSS sg13g2_decap_8
XFILLER_19_567 VDD VSS sg13g2_decap_8
XFILLER_34_504 VDD VSS sg13g2_decap_8
XFILLER_74_695 VDD VSS sg13g2_decap_8
XFILLER_73_194 VDD VSS sg13g2_decap_8
XFILLER_62_857 VDD VSS sg13g2_decap_8
XFILLER_61_312 VDD VSS sg13g2_decap_8
XFILLER_46_386 VDD VSS sg13g2_decap_8
X_1940_ _2003_/B _1940_/A _1999_/A VDD VSS sg13g2_xnor2_1
XFILLER_42_581 VDD VSS sg13g2_decap_8
XFILLER_30_721 VDD VSS sg13g2_decap_8
XFILLER_15_784 VDD VSS sg13g2_decap_8
X_1871_ VDD _2162_/A _2086_/A VSS sg13g2_inv_1
XFILLER_14_294 VDD VSS sg13g2_decap_8
XFILLER_9_77 VDD VSS sg13g2_decap_8
XFILLER_80_70 VDD VSS sg13g2_decap_8
XFILLER_31_1001 VDD VSS sg13g2_decap_8
XFILLER_30_798 VDD VSS sg13g2_decap_8
XFILLER_7_994 VDD VSS sg13g2_decap_8
X_2354_ _2354_/RESET_B VSS VDD _2354_/D _2354_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_111_553 VDD VSS sg13g2_decap_8
X_1305_ VDD _2182_/D _1305_/A VSS sg13g2_inv_1
XFILLER_96_231 VDD VSS sg13g2_decap_8
XFILLER_57_618 VDD VSS sg13g2_decap_8
XFILLER_9_1057 VDD VSS sg13g2_decap_4
XFILLER_29_0 VDD VSS sg13g2_decap_8
XFILLER_38_821 VDD VSS sg13g2_decap_8
XFILLER_56_117 VDD VSS sg13g2_decap_8
X_2285_ _2285_/RESET_B VSS VDD _2285_/D _2285_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_84_459 VDD VSS sg13g2_decap_8
XFILLER_65_651 VDD VSS sg13g2_decap_8
X_1236_ _1500_/B _1236_/C _1236_/Y VDD VSS _1226_/B sg13g2_nand3b_1
XFILLER_92_470 VDD VSS sg13g2_decap_8
XFILLER_53_824 VDD VSS sg13g2_decap_8
XFILLER_38_898 VDD VSS sg13g2_decap_8
XFILLER_64_150 VDD VSS sg13g2_decap_8
XFILLER_25_504 VDD VSS sg13g2_decap_8
XFILLER_37_364 VDD VSS sg13g2_decap_8
XFILLER_52_334 VDD VSS sg13g2_decap_8
XFILLER_52_345 VDD VSS sg13g2_fill_2
XFILLER_100_14 VDD VSS sg13g2_decap_8
XFILLER_33_581 VDD VSS sg13g2_decap_8
XFILLER_21_721 VDD VSS sg13g2_decap_8
XFILLER_52_389 VDD VSS sg13g2_fill_2
XFILLER_20_231 VDD VSS sg13g2_decap_8
XFILLER_21_798 VDD VSS sg13g2_decap_8
XFILLER_109_56 VDD VSS sg13g2_decap_8
XFILLER_106_358 VDD VSS sg13g2_decap_8
XFILLER_107_7 VDD VSS sg13g2_decap_8
XFILLER_69_49 VDD VSS sg13g2_decap_8
Xin_data_pads\[4\].in_data_pad IOVDD IOVSS _1379_/A in_data_PADs[4] VDD VSS sg13g2_IOPadIn
XFILLER_88_743 VDD VSS sg13g2_decap_8
XFILLER_88_721 VDD VSS sg13g2_decap_4
XFILLER_47_1041 VDD VSS sg13g2_decap_8
XFILLER_102_542 VDD VSS sg13g2_decap_8
XFILLER_75_404 VDD VSS sg13g2_decap_8
XFILLER_0_658 VDD VSS sg13g2_decap_8
XFILLER_87_297 VDD VSS sg13g2_fill_2
XFILLER_91_919 VDD VSS sg13g2_decap_8
XFILLER_56_651 VDD VSS sg13g2_decap_8
XFILLER_29_854 VDD VSS sg13g2_decap_8
XFILLER_18_42 VDD VSS sg13g2_decap_8
XFILLER_47_139 VDD VSS sg13g2_decap_8
XFILLER_16_504 VDD VSS sg13g2_decap_8
XFILLER_55_161 VDD VSS sg13g2_decap_8
XFILLER_28_364 VDD VSS sg13g2_decap_8
XFILLER_71_654 VDD VSS sg13g2_decap_8
XFILLER_44_879 VDD VSS sg13g2_decap_8
XFILLER_31_518 VDD VSS sg13g2_decap_8
XFILLER_70_175 VDD VSS sg13g2_decap_8
XFILLER_54_1023 VDD VSS sg13g2_fill_2
XFILLER_24_581 VDD VSS sg13g2_decap_8
XFILLER_12_721 VDD VSS sg13g2_decap_8
XFILLER_34_63 VDD VSS sg13g2_decap_8
XFILLER_43_378 VDD VSS sg13g2_decap_8
XFILLER_11_231 VDD VSS sg13g2_decap_8
XFILLER_8_714 VDD VSS sg13g2_decap_8
XFILLER_12_798 VDD VSS sg13g2_decap_8
XFILLER_15_1029 VDD VSS sg13g2_decap_8
XFILLER_7_224 VDD VSS sg13g2_decap_8
XFILLER_50_51 VDD VSS sg13g2_decap_8
XFILLER_109_196 VDD VSS sg13g2_decap_8
XFILLER_4_931 VDD VSS sg13g2_decap_8
XFILLER_98_518 VDD VSS sg13g2_decap_8
XFILLER_3_441 VDD VSS sg13g2_decap_8
XFILLER_106_881 VDD VSS sg13g2_decap_8
XFILLER_79_743 VDD VSS sg13g2_decap_8
XFILLER_61_1005 VDD VSS sg13g2_decap_8
XFILLER_22_7 VDD VSS sg13g2_decap_8
XFILLER_59_82 VDD VSS sg13g2_decap_4
XFILLER_94_713 VDD VSS sg13g2_decap_8
XFILLER_94_779 VDD VSS sg13g2_decap_8
X_2070_ _2057_/X _2069_/X _2079_/S _2071_/C VDD VSS sg13g2_mux2_1
XFILLER_93_289 VDD VSS sg13g2_decap_8
XFILLER_75_70 VDD VSS sg13g2_decap_8
XFILLER_47_684 VDD VSS sg13g2_decap_8
XFILLER_47_651 VDD VSS sg13g2_decap_8
XFILLER_19_364 VDD VSS sg13g2_decap_8
XFILLER_90_930 VDD VSS sg13g2_decap_8
XFILLER_62_610 VDD VSS sg13g2_decap_8
XFILLER_34_301 VDD VSS sg13g2_decap_8
XFILLER_90_963 VDD VSS sg13g2_fill_1
XFILLER_50_805 VDD VSS sg13g2_decap_8
XFILLER_35_868 VDD VSS sg13g2_decap_8
XFILLER_15_581 VDD VSS sg13g2_decap_8
XFILLER_61_164 VDD VSS sg13g2_decap_8
XFILLER_22_518 VDD VSS sg13g2_decap_8
XFILLER_34_378 VDD VSS sg13g2_decap_8
X_1923_ _1921_/Y _1922_/Y _1954_/S _1924_/B VDD VSS sg13g2_mux2_1
XFILLER_91_91 VDD VSS sg13g2_decap_8
XFILLER_30_595 VDD VSS sg13g2_decap_8
X_1854_ _1866_/A _1854_/C _1854_/A _1869_/A VDD VSS sg13g2_nand3_1
XIO_FILL_IO_SOUTH_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_1785_ _1900_/B _2213_/Q _2221_/Q VDD VSS sg13g2_xnor2_1
Xfanout7 _2054_/S _2021_/S VDD VSS sg13g2_buf_1
XFILLER_7_791 VDD VSS sg13g2_decap_8
XFILLER_112_840 VDD VSS sg13g2_decap_8
XFILLER_69_253 VDD VSS sg13g2_decap_8
XFILLER_97_584 VDD VSS sg13g2_decap_8
XFILLER_85_735 VDD VSS sg13g2_decap_8
X_2337_ _2337_/RESET_B VSS VDD _2337_/D _2337_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_111_350 VDD VSS sg13g2_decap_8
XFILLER_57_404 VDD VSS sg13g2_decap_8
XFILLER_73_919 VDD VSS sg13g2_fill_2
XFILLER_73_908 VDD VSS sg13g2_decap_8
XFILLER_84_234 VDD VSS sg13g2_decap_8
X_2268_ _2268_/RESET_B VSS VDD _2268_/D _2268_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_84_278 VDD VSS sg13g2_decap_8
XFILLER_72_407 VDD VSS sg13g2_decap_8
X_1219_ _1236_/C _1502_/A _2364_/D VDD VSS sg13g2_and2_1
X_2199_ _2199_/RESET_B VSS VDD _2199_/D _2199_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_66_993 VDD VSS sg13g2_decap_8
XFILLER_38_695 VDD VSS sg13g2_decap_8
XFILLER_37_161 VDD VSS sg13g2_decap_8
XFILLER_25_301 VDD VSS sg13g2_decap_8
XFILLER_81_974 VDD VSS sg13g2_decap_8
XFILLER_77_1056 VDD VSS sg13g2_decap_4
XFILLER_111_35 VDD VSS sg13g2_decap_8
XFILLER_26_868 VDD VSS sg13g2_decap_8
XFILLER_52_131 VDD VSS sg13g2_decap_8
XFILLER_80_495 VDD VSS sg13g2_decap_8
XFILLER_71_28 VDD VSS sg13g2_decap_8
XFILLER_13_518 VDD VSS sg13g2_decap_8
XFILLER_25_378 VDD VSS sg13g2_decap_8
XFILLER_21_595 VDD VSS sg13g2_decap_8
XFILLER_5_728 VDD VSS sg13g2_decap_8
XFILLER_106_133 VDD VSS sg13g2_decap_8
XFILLER_4_238 VDD VSS sg13g2_decap_8
XFILLER_20_21 VDD VSS sg13g2_decap_8
XFILLER_84_1016 VDD VSS sg13g2_decap_8
XFILLER_107_667 VDD VSS sg13g2_decap_8
XFILLER_96_14 VDD VSS sg13g2_decap_8
XFILLER_20_98 VDD VSS sg13g2_decap_8
XFILLER_1_945 VDD VSS sg13g2_decap_8
XFILLER_0_455 VDD VSS sg13g2_decap_8
XFILLER_103_884 VDD VSS sg13g2_fill_2
XFILLER_76_713 VDD VSS sg13g2_decap_8
XFILLER_102_361 VDD VSS sg13g2_decap_8
XFILLER_49_938 VDD VSS sg13g2_decap_8
XFILLER_60_1060 VDD VSS sg13g2_fill_1
XFILLER_64_908 VDD VSS sg13g2_decap_8
XFILLER_29_63 VDD VSS sg13g2_decap_8
XFILLER_48_437 VDD VSS sg13g2_decap_8
XFILLER_75_278 VDD VSS sg13g2_decap_8
XFILLER_21_1022 VDD VSS sg13g2_decap_8
XFILLER_29_651 VDD VSS sg13g2_decap_8
XFILLER_91_738 VDD VSS sg13g2_decap_8
XFILLER_57_993 VDD VSS sg13g2_decap_8
XFILLER_16_301 VDD VSS sg13g2_decap_8
XFILLER_28_161 VDD VSS sg13g2_decap_8
XFILLER_44_676 VDD VSS sg13g2_decap_8
XFILLER_44_665 VDD VSS sg13g2_fill_2
XFILLER_32_805 VDD VSS sg13g2_decap_8
XFILLER_17_868 VDD VSS sg13g2_decap_8
X_2215__110 VDD VSS _2215_/RESET_B sg13g2_tiehi
XFILLER_71_495 VDD VSS sg13g2_decap_8
XFILLER_16_378 VDD VSS sg13g2_decap_8
XFILLER_45_84 VDD VSS sg13g2_decap_8
XFILLER_31_315 VDD VSS sg13g2_decap_8
XFILLER_43_175 VDD VSS sg13g2_decap_8
XFILLER_8_511 VDD VSS sg13g2_decap_8
XFILLER_40_893 VDD VSS sg13g2_decap_8
XFILLER_12_595 VDD VSS sg13g2_decap_8
XFILLER_8_588 VDD VSS sg13g2_decap_8
X_1570_ _1577_/S0 _2241_/Q _2233_/Q _2225_/Q _2217_/Q _2287_/Q _1571_/A VDD VSS sg13g2_mux4_1
XFILLER_6_56 VDD VSS sg13g2_decap_8
XFILLER_79_540 VDD VSS sg13g2_decap_8
XFILLER_112_147 VDD VSS sg13g2_decap_8
XFILLER_79_584 VDD VSS sg13g2_decap_8
XFILLER_39_415 VDD VSS sg13g2_decap_8
XFILLER_86_91 VDD VSS sg13g2_fill_2
X_2122_ VSS VDD _2117_/Y _2120_/Y _2122_/Y _2121_/Y sg13g2_a21oi_1
XFILLER_66_223 VDD VSS sg13g2_decap_8
XFILLER_66_234 VDD VSS sg13g2_fill_1
XFILLER_94_587 VDD VSS sg13g2_decap_8
XFILLER_82_716 VDD VSS sg13g2_decap_8
XFILLER_48_960 VDD VSS sg13g2_fill_2
XFILLER_54_418 VDD VSS sg13g2_decap_8
X_2053_ _2052_/Y VDD _2336_/D VSS _2025_/A _2075_/B sg13g2_o21ai_1
XFILLER_19_161 VDD VSS sg13g2_decap_8
XFILLER_47_481 VDD VSS sg13g2_decap_8
XFILLER_63_963 VDD VSS sg13g2_fill_2
XFILLER_35_665 VDD VSS sg13g2_decap_8
XFILLER_23_805 VDD VSS sg13g2_decap_8
XFILLER_63_996 VDD VSS sg13g2_decap_8
XFILLER_62_484 VDD VSS sg13g2_decap_8
XFILLER_22_315 VDD VSS sg13g2_decap_8
XFILLER_34_175 VDD VSS sg13g2_decap_8
XFILLER_96_0 VDD VSS sg13g2_decap_8
XFILLER_50_657 VDD VSS sg13g2_decap_8
XFILLER_31_882 VDD VSS sg13g2_decap_8
X_2233__287 VDD VSS _2233_/RESET_B sg13g2_tiehi
X_1906_ _1906_/Y _1907_/A _1907_/B VDD VSS sg13g2_nand2_1
XFILLER_30_392 VDD VSS sg13g2_decap_8
X_1837_ _1921_/A _2247_/Q _2206_/Q VDD VSS sg13g2_xnor2_1
Xhold511 _2282_/Q VDD VSS hold511/X sg13g2_dlygate4sd3_1
Xhold500 _2294_/Q VDD VSS hold500/X sg13g2_dlygate4sd3_1
X_1768_ _1927_/A _1769_/B _1948_/B VDD VSS sg13g2_nor2_1
Xhold544 _1636_/Y VDD VSS _2296_/D sg13g2_dlygate4sd3_1
Xhold533 _1631_/Y VDD VSS _1632_/B sg13g2_dlygate4sd3_1
Xhold522 _2261_/Q VDD VSS hold522/X sg13g2_dlygate4sd3_1
X_1699_ _1699_/Y _1720_/A _1699_/B VDD VSS sg13g2_nand2_1
XFILLER_104_626 VDD VSS sg13g2_decap_8
Xhold566 _2366_/Q VDD VSS hold566/X sg13g2_dlygate4sd3_1
Xhold555 _2265_/Q VDD VSS hold555/X sg13g2_dlygate4sd3_1
XFILLER_106_35 VDD VSS sg13g2_decap_8
XFILLER_103_147 VDD VSS sg13g2_decap_8
XFILLER_85_510 VDD VSS sg13g2_fill_1
XFILLER_44_1033 VDD VSS sg13g2_decap_8
XFILLER_58_735 VDD VSS sg13g2_decap_8
XFILLER_100_854 VDD VSS sg13g2_decap_8
XFILLER_85_554 VDD VSS sg13g2_decap_8
XFILLER_66_28 VDD VSS sg13g2_decap_8
X_2197__146 VDD VSS _2197_/RESET_B sg13g2_tiehi
XFILLER_54_941 VDD VSS sg13g2_decap_8
XFILLER_38_481 VDD VSS sg13g2_decap_8
XFILLER_26_665 VDD VSS sg13g2_decap_8
XFILLER_14_805 VDD VSS sg13g2_decap_8
XFILLER_81_793 VDD VSS sg13g2_fill_1
XFILLER_82_49 VDD VSS sg13g2_decap_8
XFILLER_53_484 VDD VSS sg13g2_decap_8
XFILLER_13_315 VDD VSS sg13g2_decap_8
XFILLER_15_21 VDD VSS sg13g2_decap_8
XFILLER_25_175 VDD VSS sg13g2_decap_8
XFILLER_41_657 VDD VSS sg13g2_decap_8
XFILLER_40_112 VDD VSS sg13g2_decap_8
XFILLER_9_308 VDD VSS sg13g2_decap_8
XFILLER_15_98 VDD VSS sg13g2_decap_8
X_2349__105 VDD VSS _2349_/RESET_B sg13g2_tiehi
XFILLER_22_882 VDD VSS sg13g2_decap_8
XFILLER_40_189 VDD VSS sg13g2_decap_8
XFILLER_51_1059 VDD VSS sg13g2_fill_2
XFILLER_31_42 VDD VSS sg13g2_decap_8
XFILLER_21_392 VDD VSS sg13g2_decap_8
X_2249__250 VDD VSS _2249_/RESET_B sg13g2_tiehi
XFILLER_5_525 VDD VSS sg13g2_decap_8
XFILLER_108_976 VDD VSS sg13g2_decap_8
XFILLER_96_808 VDD VSS sg13g2_decap_8
XFILLER_1_742 VDD VSS sg13g2_decap_8
XFILLER_95_307 VDD VSS sg13g2_decap_8
XFILLER_0_252 VDD VSS sg13g2_decap_8
XFILLER_48_267 VDD VSS sg13g2_decap_8
XFILLER_91_535 VDD VSS sg13g2_decap_8
XFILLER_56_83 VDD VSS sg13g2_decap_4
XFILLER_60_900 VDD VSS sg13g2_decap_8
XFILLER_63_248 VDD VSS sg13g2_decap_8
XFILLER_17_665 VDD VSS sg13g2_decap_8
XFILLER_45_996 VDD VSS sg13g2_decap_8
XFILLER_32_602 VDD VSS sg13g2_decap_8
XFILLER_16_175 VDD VSS sg13g2_decap_8
X_2291__145 VDD VSS _2291_/RESET_B sg13g2_tiehi
XFILLER_31_112 VDD VSS sg13g2_decap_8
XFILLER_44_495 VDD VSS sg13g2_decap_4
XFILLER_32_679 VDD VSS sg13g2_decap_8
XFILLER_20_819 VDD VSS sg13g2_decap_8
XFILLER_40_690 VDD VSS sg13g2_decap_8
XFILLER_13_882 VDD VSS sg13g2_decap_8
XFILLER_31_189 VDD VSS sg13g2_decap_8
XFILLER_12_392 VDD VSS sg13g2_decap_8
XFILLER_9_875 VDD VSS sg13g2_decap_8
XFILLER_8_385 VDD VSS sg13g2_decap_8
X_1622_ _1628_/A _2294_/Q _2279_/Q VDD VSS sg13g2_xnor2_1
XFILLER_99_646 VDD VSS sg13g2_fill_2
XFILLER_98_112 VDD VSS sg13g2_decap_8
X_1553_ _1552_/Y VDD _1553_/Y VSS _1592_/A _1550_/Y sg13g2_o21ai_1
XFILLER_87_808 VDD VSS sg13g2_decap_8
X_1484_ _2364_/Q _2355_/Q _1487_/B VDD VSS sg13g2_nor2_1
XFILLER_101_629 VDD VSS sg13g2_decap_8
XFILLER_79_370 VDD VSS sg13g2_decap_8
XFILLER_67_532 VDD VSS sg13g2_decap_8
XFILLER_11_0 VDD VSS sg13g2_decap_8
XFILLER_39_245 VDD VSS sg13g2_decap_8
XFILLER_95_896 VDD VSS sg13g2_decap_8
XFILLER_94_384 VDD VSS sg13g2_decap_8
XFILLER_82_513 VDD VSS sg13g2_decap_8
XFILLER_55_727 VDD VSS sg13g2_decap_8
X_2105_ VSS VDD _2102_/B _2102_/C _2105_/Y _2102_/A sg13g2_a21oi_1
X_2036_ _2026_/X _1826_/B _2036_/S _2037_/B VDD VSS sg13g2_mux2_1
XFILLER_36_952 VDD VSS sg13g2_decap_8
XFILLER_63_793 VDD VSS sg13g2_decap_8
XFILLER_51_911 VDD VSS sg13g2_decap_8
XFILLER_23_602 VDD VSS sg13g2_decap_8
XFILLER_35_462 VDD VSS sg13g2_decap_8
XFILLER_74_1059 VDD VSS sg13g2_fill_2
XFILLER_22_112 VDD VSS sg13g2_decap_8
XFILLER_23_679 VDD VSS sg13g2_decap_8
XFILLER_11_819 VDD VSS sg13g2_decap_8
XFILLER_50_465 VDD VSS sg13g2_decap_8
XFILLER_10_329 VDD VSS sg13g2_decap_8
XFILLER_22_189 VDD VSS sg13g2_decap_8
XFILLER_109_707 VDD VSS sg13g2_decap_8
XFILLER_11_1043 VDD VSS sg13g2_decap_8
XFILLER_105_924 VDD VSS sg13g2_decap_8
Xhold352 _1294_/Y VDD VSS _1295_/A sg13g2_dlygate4sd3_1
XFILLER_89_112 VDD VSS sg13g2_decap_8
Xhold341 _1487_/Y VDD VSS hold341/X sg13g2_dlygate4sd3_1
Xhold330 _2105_/Y VDD VSS _2106_/C sg13g2_dlygate4sd3_1
XFILLER_2_539 VDD VSS sg13g2_decap_8
XFILLER_81_1008 VDD VSS sg13g2_decap_8
Xhold385 _2184_/Q VDD VSS hold385/X sg13g2_dlygate4sd3_1
Xhold363 _1326_/Y VDD VSS _1327_/A sg13g2_dlygate4sd3_1
Xhold396 _2359_/Q VDD VSS _1501_/A sg13g2_dlygate4sd3_1
Xhold374 _1473_/Y VDD VSS _2255_/D sg13g2_dlygate4sd3_1
XFILLER_77_329 VDD VSS sg13g2_decap_8
XFILLER_77_49 VDD VSS sg13g2_decap_8
XFILLER_86_830 VDD VSS sg13g2_decap_8
XFILLER_58_532 VDD VSS sg13g2_decap_4
XFILLER_100_651 VDD VSS sg13g2_fill_1
XFILLER_85_362 VDD VSS sg13g2_decap_8
XFILLER_73_524 VDD VSS sg13g2_decap_8
XFILLER_27_952 VDD VSS sg13g2_decap_8
XFILLER_26_42 VDD VSS sg13g2_decap_8
XFILLER_60_207 VDD VSS sg13g2_decap_8
XFILLER_14_602 VDD VSS sg13g2_decap_8
XFILLER_26_462 VDD VSS sg13g2_decap_8
XFILLER_42_966 VDD VSS sg13g2_decap_8
XFILLER_53_292 VDD VSS sg13g2_decap_8
XFILLER_13_112 VDD VSS sg13g2_decap_8
XFILLER_9_105 VDD VSS sg13g2_decap_8
XFILLER_14_679 VDD VSS sg13g2_decap_8
XFILLER_41_465 VDD VSS sg13g2_fill_2
XFILLER_13_189 VDD VSS sg13g2_decap_8
XFILLER_6_812 VDD VSS sg13g2_decap_8
XFILLER_42_63 VDD VSS sg13g2_decap_8
XFILLER_5_322 VDD VSS sg13g2_decap_8
XFILLER_10_896 VDD VSS sg13g2_decap_8
XFILLER_108_773 VDD VSS sg13g2_decap_8
XFILLER_6_889 VDD VSS sg13g2_decap_8
XFILLER_5_399 VDD VSS sg13g2_decap_8
XFILLER_111_938 VDD VSS sg13g2_decap_8
XFILLER_96_616 VDD VSS sg13g2_decap_8
XFILLER_3_35 VDD VSS sg13g2_decap_8
XFILLER_77_830 VDD VSS sg13g2_decap_8
XFILLER_95_126 VDD VSS sg13g2_decap_8
XFILLER_27_1050 VDD VSS sg13g2_decap_8
XFILLER_49_521 VDD VSS sg13g2_decap_4
XFILLER_77_863 VDD VSS sg13g2_decap_8
XFILLER_110_459 VDD VSS sg13g2_decap_8
XFILLER_76_340 VDD VSS sg13g2_fill_1
XFILLER_49_565 VDD VSS sg13g2_decap_8
XFILLER_3_1008 VDD VSS sg13g2_decap_8
XFILLER_92_833 VDD VSS sg13g2_decap_8
XFILLER_76_373 VDD VSS sg13g2_decap_8
XFILLER_37_749 VDD VSS sg13g2_decap_8
XFILLER_64_557 VDD VSS sg13g2_decap_8
XFILLER_18_952 VDD VSS sg13g2_decap_8
XFILLER_36_259 VDD VSS sg13g2_decap_8
XFILLER_92_899 VDD VSS sg13g2_decap_8
XFILLER_83_70 VDD VSS sg13g2_decap_8
XFILLER_52_719 VDD VSS sg13g2_decap_8
XFILLER_17_462 VDD VSS sg13g2_decap_8
XFILLER_33_966 VDD VSS sg13g2_decap_8
XFILLER_20_616 VDD VSS sg13g2_decap_8
XFILLER_34_1043 VDD VSS sg13g2_decap_8
XFILLER_60_785 VDD VSS sg13g2_decap_8
XFILLER_32_476 VDD VSS sg13g2_decap_8
XFILLER_9_672 VDD VSS sg13g2_decap_8
XFILLER_8_182 VDD VSS sg13g2_decap_8
XFILLER_59_0 VDD VSS sg13g2_decap_8
X_1605_ _1606_/B _2291_/Q _2276_/Q VDD VSS sg13g2_xnor2_1
X_1536_ VDD _1536_/Y _1536_/A VSS sg13g2_inv_1
XFILLER_102_916 VDD VSS sg13g2_decap_4
XFILLER_87_616 VDD VSS sg13g2_decap_8
XFILLER_99_476 VDD VSS sg13g2_decap_8
XFILLER_59_307 VDD VSS sg13g2_fill_1
XFILLER_102_949 VDD VSS sg13g2_decap_8
XFILLER_101_437 VDD VSS sg13g2_decap_8
XFILLER_68_841 VDD VSS sg13g2_decap_8
X_1467_ VSS VDD _1201_/Y _1481_/A2 _2252_/D _1466_/Y sg13g2_a21oi_1
X_1398_ VDD _2221_/D _1398_/A VSS sg13g2_inv_1
XFILLER_41_1014 VDD VSS sg13g2_decap_8
XFILLER_95_693 VDD VSS sg13g2_decap_8
XFILLER_83_822 VDD VSS sg13g2_decap_8
XFILLER_103_14 VDD VSS sg13g2_decap_8
XFILLER_28_749 VDD VSS sg13g2_decap_8
XFILLER_82_321 VDD VSS sg13g2_decap_8
XFILLER_55_546 VDD VSS sg13g2_decap_8
XFILLER_27_259 VDD VSS sg13g2_decap_8
XFILLER_83_899 VDD VSS sg13g2_decap_8
XFILLER_82_387 VDD VSS sg13g2_decap_8
XFILLER_70_505 VDD VSS sg13g2_decap_8
XFILLER_70_516 VDD VSS sg13g2_fill_1
X_2019_ _1998_/X _2008_/X _2022_/S _2019_/X VDD VSS sg13g2_mux2_1
XFILLER_70_549 VDD VSS sg13g2_decap_8
XFILLER_51_730 VDD VSS sg13g2_fill_2
XFILLER_24_966 VDD VSS sg13g2_decap_8
XFILLER_11_616 VDD VSS sg13g2_decap_8
XFILLER_23_476 VDD VSS sg13g2_decap_8
XFILLER_109_504 VDD VSS sg13g2_decap_8
XFILLER_10_126 VDD VSS sg13g2_decap_8
XFILLER_7_609 VDD VSS sg13g2_decap_8
XFILLER_6_119 VDD VSS sg13g2_decap_8
X_2346__119 VDD VSS _2346_/RESET_B sg13g2_tiehi
XFILLER_12_77 VDD VSS sg13g2_decap_8
XFILLER_105_721 VDD VSS sg13g2_decap_8
XFILLER_3_826 VDD VSS sg13g2_decap_8
XFILLER_104_231 VDD VSS sg13g2_decap_8
X_2246__253 VDD VSS _2246_/RESET_B sg13g2_tiehi
XFILLER_2_336 VDD VSS sg13g2_decap_8
XFILLER_105_798 VDD VSS sg13g2_decap_8
XFILLER_77_126 VDD VSS sg13g2_decap_8
XFILLER_74_800 VDD VSS sg13g2_decap_8
XFILLER_58_351 VDD VSS sg13g2_decap_8
XFILLER_86_693 VDD VSS sg13g2_decap_8
XFILLER_19_749 VDD VSS sg13g2_decap_8
XFILLER_46_524 VDD VSS sg13g2_decap_8
XFILLER_85_192 VDD VSS sg13g2_decap_8
XFILLER_18_259 VDD VSS sg13g2_decap_8
XFILLER_37_63 VDD VSS sg13g2_decap_8
XFILLER_73_365 VDD VSS sg13g2_decap_8
XFILLER_57_1010 VDD VSS sg13g2_decap_8
XFILLER_61_505 VDD VSS sg13g2_decap_4
XFILLER_42_763 VDD VSS sg13g2_decap_8
XFILLER_30_903 VDD VSS sg13g2_decap_8
XFILLER_15_966 VDD VSS sg13g2_decap_8
XFILLER_53_62 VDD VSS sg13g2_decap_8
XFILLER_105_1008 VDD VSS sg13g2_decap_8
XFILLER_14_476 VDD VSS sg13g2_decap_8
XFILLER_41_262 VDD VSS sg13g2_decap_8
X_2227__86 VDD VSS _2227__86/L_HI sg13g2_tiehi
XFILLER_10_693 VDD VSS sg13g2_decap_8
XFILLER_108_570 VDD VSS sg13g2_decap_8
XFILLER_6_686 VDD VSS sg13g2_decap_8
XFILLER_52_7 VDD VSS sg13g2_decap_8
XFILLER_64_1014 VDD VSS sg13g2_decap_8
XFILLER_5_196 VDD VSS sg13g2_decap_8
X_2370_ _2370__85/L_HI VSS VDD _2370_/D _2370_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_96_413 VDD VSS sg13g2_decap_8
XFILLER_111_735 VDD VSS sg13g2_decap_8
X_1321_ VDD _2190_/D _1321_/A VSS sg13g2_inv_1
XFILLER_69_649 VDD VSS sg13g2_decap_8
XFILLER_78_70 VDD VSS sg13g2_decap_8
XFILLER_77_660 VDD VSS sg13g2_decap_8
XFILLER_110_245 VDD VSS sg13g2_decap_8
XFILLER_96_479 VDD VSS sg13g2_decap_8
X_1252_ _1252_/Y _1252_/B _1250_/B VDD VSS sg13g2_nand2b_1
XFILLER_49_351 VDD VSS sg13g2_fill_2
XFILLER_49_384 VDD VSS sg13g2_decap_8
XFILLER_37_546 VDD VSS sg13g2_decap_8
XFILLER_64_321 VDD VSS sg13g2_decap_8
XFILLER_80_825 VDD VSS sg13g2_decap_8
XFILLER_94_91 VDD VSS sg13g2_decap_8
XFILLER_65_888 VDD VSS sg13g2_decap_8
XFILLER_52_505 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_92_696 VDD VSS sg13g2_decap_8
XFILLER_33_763 VDD VSS sg13g2_decap_8
XFILLER_21_903 VDD VSS sg13g2_decap_8
XFILLER_20_413 VDD VSS sg13g2_decap_8
XFILLER_32_273 VDD VSS sg13g2_decap_8
XFILLER_106_518 VDD VSS sg13g2_decap_8
XFILLER_88_914 VDD VSS sg13g2_decap_8
XFILLER_87_402 VDD VSS sg13g2_decap_8
X_1519_ VSS VDD _2120_/A hold546/X _2273_/D _1261_/Y sg13g2_a21oi_1
XFILLER_101_234 VDD VSS sg13g2_decap_8
XFILLER_87_468 VDD VSS sg13g2_decap_8
XFILLER_95_490 VDD VSS sg13g2_decap_4
XFILLER_74_28 VDD VSS sg13g2_decap_8
XFILLER_28_546 VDD VSS sg13g2_decap_8
XFILLER_67_181 VDD VSS sg13g2_decap_8
XFILLER_55_343 VDD VSS sg13g2_fill_1
XFILLER_83_663 VDD VSS sg13g2_decap_8
XFILLER_56_899 VDD VSS sg13g2_decap_8
XFILLER_43_516 VDD VSS sg13g2_fill_1
XFILLER_43_505 VDD VSS sg13g2_decap_8
XFILLER_71_847 VDD VSS sg13g2_decap_8
XFILLER_70_313 VDD VSS sg13g2_decap_8
XFILLER_70_379 VDD VSS sg13g2_decap_8
XFILLER_24_763 VDD VSS sg13g2_decap_8
XFILLER_12_903 VDD VSS sg13g2_decap_8
XFILLER_90_49 VDD VSS sg13g2_decap_8
XFILLER_11_413 VDD VSS sg13g2_decap_8
XFILLER_23_21 VDD VSS sg13g2_decap_8
XFILLER_23_273 VDD VSS sg13g2_decap_8
XFILLER_51_593 VDD VSS sg13g2_decap_8
XFILLER_7_406 VDD VSS sg13g2_decap_8
XFILLER_104_1041 VDD VSS sg13g2_decap_8
XFILLER_20_980 VDD VSS sg13g2_decap_8
XFILLER_99_14 VDD VSS sg13g2_decap_8
XFILLER_23_98 VDD VSS sg13g2_decap_8
XFILLER_87_1047 VDD VSS sg13g2_decap_8
XFILLER_48_1009 VDD VSS sg13g2_decap_8
XFILLER_3_623 VDD VSS sg13g2_decap_8
XFILLER_105_540 VDD VSS sg13g2_decap_8
XFILLER_2_133 VDD VSS sg13g2_decap_8
XFILLER_79_947 VDD VSS sg13g2_decap_8
XFILLER_105_595 VDD VSS sg13g2_decap_8
XFILLER_78_424 VDD VSS sg13g2_fill_2
XFILLER_94_906 VDD VSS sg13g2_decap_8
XFILLER_78_468 VDD VSS sg13g2_decap_8
XFILLER_111_1001 VDD VSS sg13g2_decap_8
XFILLER_59_671 VDD VSS sg13g2_decap_8
XFILLER_93_449 VDD VSS sg13g2_decap_8
XFILLER_47_866 VDD VSS sg13g2_decap_8
XFILLER_0_14 VDD VSS sg13g2_decap_8
XFILLER_19_546 VDD VSS sg13g2_decap_8
XFILLER_94_1018 VDD VSS sg13g2_decap_8
XFILLER_74_674 VDD VSS sg13g2_decap_8
XFILLER_94_1029 VDD VSS sg13g2_fill_1
XFILLER_62_836 VDD VSS sg13g2_decap_8
XFILLER_15_763 VDD VSS sg13g2_decap_8
XFILLER_30_700 VDD VSS sg13g2_decap_8
XFILLER_14_273 VDD VSS sg13g2_decap_8
X_1870_ _1870_/B _1870_/A _2086_/A VDD VSS sg13g2_xor2_1
XFILLER_9_56 VDD VSS sg13g2_decap_8
XFILLER_70_1051 VDD VSS sg13g2_decap_8
XFILLER_30_777 VDD VSS sg13g2_decap_8
XFILLER_31_1057 VDD VSS sg13g2_decap_4
XFILLER_11_980 VDD VSS sg13g2_decap_8
XFILLER_10_490 VDD VSS sg13g2_decap_8
XFILLER_7_973 VDD VSS sg13g2_decap_8
XFILLER_6_483 VDD VSS sg13g2_decap_8
XFILLER_89_91 VDD VSS sg13g2_decap_8
XFILLER_97_733 VDD VSS sg13g2_fill_1
XFILLER_97_722 VDD VSS sg13g2_decap_8
XFILLER_96_210 VDD VSS sg13g2_decap_8
X_2353_ _2353_/RESET_B VSS VDD _2353_/D _2353_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_9_1036 VDD VSS sg13g2_decap_8
X_1304_ _1304_/Y _1322_/B1 hold364/X _1322_/A2 _2346_/Q VDD VSS sg13g2_a22oi_1
XFILLER_111_532 VDD VSS sg13g2_decap_8
XFILLER_96_287 VDD VSS sg13g2_decap_8
XFILLER_38_800 VDD VSS sg13g2_decap_8
X_2284_ _2284_/RESET_B VSS VDD _2284_/D _2284_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_65_641 VDD VSS sg13g2_decap_4
X_1235_ _1235_/A _1409_/C _2261_/D VDD VSS sg13g2_nor2_1
XFILLER_93_972 VDD VSS sg13g2_decap_8
XFILLER_38_877 VDD VSS sg13g2_decap_8
XFILLER_37_343 VDD VSS sg13g2_decap_8
XFILLER_80_644 VDD VSS sg13g2_decap_4
XFILLER_65_696 VDD VSS sg13g2_decap_8
XFILLER_52_368 VDD VSS sg13g2_decap_8
XFILLER_33_560 VDD VSS sg13g2_decap_8
XFILLER_21_700 VDD VSS sg13g2_decap_8
XFILLER_40_519 VDD VSS sg13g2_decap_8
XFILLER_20_210 VDD VSS sg13g2_decap_8
XFILLER_21_777 VDD VSS sg13g2_decap_8
X_1999_ _2022_/S _2021_/S _1999_/A _2033_/B VDD VSS sg13g2_nand3_1
XFILLER_20_287 VDD VSS sg13g2_decap_8
XFILLER_109_35 VDD VSS sg13g2_decap_8
XFILLER_107_849 VDD VSS sg13g2_decap_8
XFILLER_106_326 VDD VSS sg13g2_decap_8
XFILLER_69_28 VDD VSS sg13g2_decap_8
XFILLER_88_700 VDD VSS sg13g2_decap_8
XFILLER_47_1020 VDD VSS sg13g2_decap_8
XFILLER_102_521 VDD VSS sg13g2_decap_8
X_2243__256 VDD VSS _2243_/RESET_B sg13g2_tiehi
XFILLER_0_637 VDD VSS sg13g2_decap_8
XFILLER_88_788 VDD VSS sg13g2_decap_8
XFILLER_87_276 VDD VSS sg13g2_decap_8
XFILLER_85_49 VDD VSS sg13g2_decap_8
XFILLER_75_449 VDD VSS sg13g2_fill_1
XFILLER_56_630 VDD VSS sg13g2_decap_8
XFILLER_29_833 VDD VSS sg13g2_decap_8
XFILLER_18_21 VDD VSS sg13g2_decap_8
XFILLER_84_961 VDD VSS sg13g2_decap_4
XFILLER_44_825 VDD VSS sg13g2_decap_8
XFILLER_55_140 VDD VSS sg13g2_decap_8
XFILLER_28_343 VDD VSS sg13g2_decap_8
XFILLER_84_994 VDD VSS sg13g2_decap_8
XFILLER_71_633 VDD VSS sg13g2_decap_8
XFILLER_44_858 VDD VSS sg13g2_decap_8
XFILLER_44_836 VDD VSS sg13g2_fill_2
XFILLER_18_98 VDD VSS sg13g2_decap_8
XFILLER_70_154 VDD VSS sg13g2_decap_8
XFILLER_43_357 VDD VSS sg13g2_decap_8
XFILLER_71_699 VDD VSS sg13g2_decap_8
XFILLER_24_560 VDD VSS sg13g2_decap_8
XFILLER_12_700 VDD VSS sg13g2_decap_8
XFILLER_34_42 VDD VSS sg13g2_decap_8
XFILLER_54_1057 VDD VSS sg13g2_decap_4
X_2250__249 VDD VSS _2250_/RESET_B sg13g2_tiehi
XFILLER_11_210 VDD VSS sg13g2_decap_8
XFILLER_15_1008 VDD VSS sg13g2_decap_8
XFILLER_7_203 VDD VSS sg13g2_decap_8
XFILLER_12_777 VDD VSS sg13g2_decap_8
XFILLER_11_287 VDD VSS sg13g2_decap_8
XFILLER_50_30 VDD VSS sg13g2_fill_1
XFILLER_4_910 VDD VSS sg13g2_decap_8
X_2287__161 VDD VSS _2287_/RESET_B sg13g2_tiehi
XFILLER_109_175 VDD VSS sg13g2_decap_8
XFILLER_3_420 VDD VSS sg13g2_decap_8
XFILLER_106_860 VDD VSS sg13g2_decap_8
XFILLER_4_987 VDD VSS sg13g2_decap_8
XFILLER_79_722 VDD VSS sg13g2_decap_8
XFILLER_112_329 VDD VSS sg13g2_decap_8
XFILLER_3_497 VDD VSS sg13g2_decap_8
XFILLER_67_917 VDD VSS sg13g2_decap_4
XFILLER_93_213 VDD VSS sg13g2_decap_8
XFILLER_39_619 VDD VSS sg13g2_decap_8
XFILLER_93_235 VDD VSS sg13g2_fill_1
XFILLER_47_630 VDD VSS sg13g2_decap_8
XFILLER_66_449 VDD VSS sg13g2_decap_8
XFILLER_59_490 VDD VSS sg13g2_decap_8
XFILLER_15_7 VDD VSS sg13g2_decap_8
XFILLER_93_257 VDD VSS sg13g2_decap_8
XFILLER_81_419 VDD VSS sg13g2_decap_8
XFILLER_19_343 VDD VSS sg13g2_decap_8
XFILLER_74_493 VDD VSS sg13g2_decap_8
XFILLER_35_847 VDD VSS sg13g2_decap_8
XFILLER_62_655 VDD VSS sg13g2_decap_8
XFILLER_61_143 VDD VSS sg13g2_decap_8
XFILLER_34_357 VDD VSS sg13g2_decap_8
XFILLER_15_560 VDD VSS sg13g2_decap_8
X_1922_ VSS VDD _1906_/Y _1921_/Y _1922_/Y _1952_/B sg13g2_a21oi_1
XFILLER_91_70 VDD VSS sg13g2_decap_8
XFILLER_43_891 VDD VSS sg13g2_decap_8
XFILLER_30_574 VDD VSS sg13g2_decap_8
X_1853_ _1854_/C _2251_/Q _2210_/Q VDD VSS sg13g2_xnor2_1
XIO_BOND_in_data_pads\[3\].in_data_pad in_data_PADs[3] bondpad_70x70
X_1784_ _1780_/Y VDD _1900_/A VSS _1929_/A _1782_/Y sg13g2_o21ai_1
XFILLER_7_770 VDD VSS sg13g2_decap_8
Xfanout8 _1997_/Y _2054_/S VDD VSS sg13g2_buf_1
XFILLER_6_280 VDD VSS sg13g2_decap_8
XFILLER_89_508 VDD VSS sg13g2_decap_8
XFILLER_41_0 VDD VSS sg13g2_decap_8
XFILLER_97_530 VDD VSS sg13g2_decap_8
XFILLER_112_896 VDD VSS sg13g2_decap_8
XFILLER_97_563 VDD VSS sg13g2_decap_8
XFILLER_85_703 VDD VSS sg13g2_fill_1
XFILLER_84_202 VDD VSS sg13g2_fill_1
X_2336_ _2336_/RESET_B VSS VDD _2336_/D _2336_/Q clkload8/A sg13g2_dfrbpq_1
X_2267_ _2267_/RESET_B VSS VDD _2267_/D _2267_/Q _2289_/CLK sg13g2_dfrbpq_1
X_1218_ VDD _1218_/Y _2243_/Q VSS sg13g2_inv_1
XFILLER_38_674 VDD VSS sg13g2_decap_8
XFILLER_37_140 VDD VSS sg13g2_decap_8
XFILLER_77_1035 VDD VSS sg13g2_decap_8
XFILLER_93_780 VDD VSS sg13g2_decap_8
X_2198_ _2198_/RESET_B VSS VDD _2198_/D _2198_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_26_847 VDD VSS sg13g2_decap_8
XFILLER_52_110 VDD VSS sg13g2_decap_8
XFILLER_81_953 VDD VSS sg13g2_decap_8
XFILLER_111_14 VDD VSS sg13g2_decap_8
XFILLER_53_666 VDD VSS sg13g2_decap_8
XFILLER_25_357 VDD VSS sg13g2_decap_8
XFILLER_80_474 VDD VSS sg13g2_decap_8
XFILLER_53_677 VDD VSS sg13g2_fill_1
XFILLER_41_839 VDD VSS sg13g2_decap_8
XFILLER_40_349 VDD VSS sg13g2_decap_8
XFILLER_21_574 VDD VSS sg13g2_decap_8
XFILLER_5_707 VDD VSS sg13g2_decap_8
XFILLER_101_1055 VDD VSS sg13g2_decap_4
XFILLER_107_646 VDD VSS sg13g2_decap_8
XFILLER_106_112 VDD VSS sg13g2_decap_8
XFILLER_4_217 VDD VSS sg13g2_decap_8
XFILLER_20_77 VDD VSS sg13g2_decap_8
XFILLER_106_189 VDD VSS sg13g2_decap_8
XFILLER_1_924 VDD VSS sg13g2_decap_8
XFILLER_88_541 VDD VSS sg13g2_fill_2
XFILLER_0_434 VDD VSS sg13g2_decap_8
XFILLER_103_896 VDD VSS sg13g2_decap_8
XFILLER_29_42 VDD VSS sg13g2_decap_8
XFILLER_48_416 VDD VSS sg13g2_decap_8
XFILLER_76_769 VDD VSS sg13g2_decap_8
XFILLER_21_1001 VDD VSS sg13g2_decap_8
XFILLER_29_630 VDD VSS sg13g2_decap_8
XFILLER_75_257 VDD VSS sg13g2_decap_8
XFILLER_63_419 VDD VSS sg13g2_fill_2
XFILLER_63_408 VDD VSS sg13g2_decap_8
XFILLER_28_140 VDD VSS sg13g2_decap_8
XFILLER_17_847 VDD VSS sg13g2_decap_8
XFILLER_90_249 VDD VSS sg13g2_decap_8
XFILLER_16_357 VDD VSS sg13g2_decap_8
XFILLER_45_63 VDD VSS sg13g2_decap_8
XFILLER_72_997 VDD VSS sg13g2_decap_8
XFILLER_71_474 VDD VSS sg13g2_decap_8
XFILLER_43_154 VDD VSS sg13g2_fill_2
XFILLER_101_91 VDD VSS sg13g2_decap_8
XFILLER_40_872 VDD VSS sg13g2_decap_8
XFILLER_12_574 VDD VSS sg13g2_decap_8
XFILLER_8_567 VDD VSS sg13g2_decap_8
XFILLER_6_35 VDD VSS sg13g2_decap_8
XFILLER_4_784 VDD VSS sg13g2_decap_8
XFILLER_112_126 VDD VSS sg13g2_decap_8
XFILLER_3_294 VDD VSS sg13g2_decap_8
XFILLER_66_202 VDD VSS sg13g2_decap_8
XFILLER_94_522 VDD VSS sg13g2_decap_8
XFILLER_86_70 VDD VSS sg13g2_decap_8
X_2121_ _1688_/B VDD _2121_/Y VSS _1259_/A hold567/X sg13g2_o21ai_1
XFILLER_67_769 VDD VSS sg13g2_decap_8
XFILLER_55_909 VDD VSS sg13g2_decap_8
X_2052_ _2052_/Y _2149_/A _2077_/A VDD VSS sg13g2_nand2_1
XFILLER_19_140 VDD VSS sg13g2_decap_8
XFILLER_81_249 VDD VSS sg13g2_decap_8
XFILLER_35_644 VDD VSS sg13g2_decap_8
XFILLER_90_794 VDD VSS sg13g2_fill_1
XFILLER_62_463 VDD VSS sg13g2_decap_8
XFILLER_34_154 VDD VSS sg13g2_decap_8
XFILLER_50_636 VDD VSS sg13g2_decap_8
XFILLER_89_0 VDD VSS sg13g2_decap_8
XFILLER_31_861 VDD VSS sg13g2_decap_8
X_1905_ _1907_/B _1905_/A _1905_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_371 VDD VSS sg13g2_decap_8
X_1836_ _1844_/B _2247_/Q _2206_/Q VDD VSS sg13g2_nand2b_1
X_1767_ _1769_/B _1926_/B _1767_/B _1940_/A VDD VSS sg13g2_and3_1
Xhold501 _1625_/Y VDD VSS _1626_/B sg13g2_dlygate4sd3_1
XFILLER_104_605 VDD VSS sg13g2_decap_8
Xhold545 _2365_/Q VDD VSS _1500_/A sg13g2_dlygate4sd3_1
Xhold512 _1582_/Y VDD VSS _1583_/B sg13g2_dlygate4sd3_1
Xhold534 _1632_/Y VDD VSS _2295_/D sg13g2_dlygate4sd3_1
Xhold523 _2291_/Q VDD VSS hold523/X sg13g2_dlygate4sd3_1
X_1698_ _1699_/B _1698_/A _1703_/A VDD VSS sg13g2_xnor2_1
Xhold567 _2367_/Q VDD VSS hold567/X sg13g2_dlygate4sd3_1
Xhold556 _1490_/Y VDD VSS _1491_/C sg13g2_dlygate4sd3_1
XFILLER_89_349 VDD VSS sg13g2_decap_8
XFILLER_106_14 VDD VSS sg13g2_decap_8
XFILLER_103_126 VDD VSS sg13g2_decap_8
XFILLER_44_1012 VDD VSS sg13g2_decap_8
XFILLER_100_800 VDD VSS sg13g2_decap_4
XFILLER_58_714 VDD VSS sg13g2_decap_8
X_2319_ _2319_/RESET_B VSS VDD _2319_/D _2319_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_112_693 VDD VSS sg13g2_decap_8
XFILLER_100_833 VDD VSS sg13g2_decap_8
XFILLER_97_393 VDD VSS sg13g2_decap_8
XFILLER_85_533 VDD VSS sg13g2_decap_8
XFILLER_57_257 VDD VSS sg13g2_fill_1
XFILLER_57_246 VDD VSS sg13g2_decap_8
XFILLER_39_983 VDD VSS sg13g2_decap_8
XFILLER_38_460 VDD VSS sg13g2_decap_8
XFILLER_81_750 VDD VSS sg13g2_decap_4
XFILLER_82_28 VDD VSS sg13g2_decap_8
XFILLER_26_644 VDD VSS sg13g2_decap_8
XFILLER_81_761 VDD VSS sg13g2_fill_1
XFILLER_54_997 VDD VSS sg13g2_decap_8
XFILLER_53_463 VDD VSS sg13g2_decap_8
XFILLER_25_154 VDD VSS sg13g2_decap_8
XFILLER_41_636 VDD VSS sg13g2_decap_8
XFILLER_90_1043 VDD VSS sg13g2_decap_8
XFILLER_22_861 VDD VSS sg13g2_decap_8
XFILLER_15_77 VDD VSS sg13g2_decap_8
XFILLER_40_168 VDD VSS sg13g2_decap_8
XFILLER_51_1038 VDD VSS sg13g2_decap_8
XFILLER_21_371 VDD VSS sg13g2_decap_8
XFILLER_5_504 VDD VSS sg13g2_decap_8
XFILLER_31_21 VDD VSS sg13g2_decap_8
XFILLER_108_955 VDD VSS sg13g2_decap_8
XFILLER_107_465 VDD VSS sg13g2_decap_8
XFILLER_31_98 VDD VSS sg13g2_decap_8
XFILLER_107_487 VDD VSS sg13g2_decap_8
XFILLER_1_721 VDD VSS sg13g2_decap_8
XFILLER_89_894 VDD VSS sg13g2_decap_8
XFILLER_0_231 VDD VSS sg13g2_decap_8
XFILLER_76_533 VDD VSS sg13g2_decap_8
XFILLER_1_798 VDD VSS sg13g2_decap_8
XFILLER_49_769 VDD VSS sg13g2_decap_8
XFILLER_5_1050 VDD VSS sg13g2_decap_8
XFILLER_91_514 VDD VSS sg13g2_decap_8
XFILLER_64_739 VDD VSS sg13g2_decap_8
XFILLER_56_51 VDD VSS sg13g2_decap_8
XFILLER_56_62 VDD VSS sg13g2_fill_1
XFILLER_17_644 VDD VSS sg13g2_decap_8
XFILLER_45_975 VDD VSS sg13g2_decap_8
XFILLER_16_154 VDD VSS sg13g2_decap_8
XFILLER_44_474 VDD VSS sg13g2_fill_2
XFILLER_72_794 VDD VSS sg13g2_decap_8
XFILLER_60_956 VDD VSS sg13g2_decap_8
XFILLER_32_658 VDD VSS sg13g2_decap_8
XFILLER_108_1039 VDD VSS sg13g2_decap_8
XFILLER_13_861 VDD VSS sg13g2_decap_8
XFILLER_31_168 VDD VSS sg13g2_decap_8
XFILLER_82_7 VDD VSS sg13g2_decap_8
XFILLER_12_371 VDD VSS sg13g2_decap_8
XFILLER_9_854 VDD VSS sg13g2_decap_8
XFILLER_8_364 VDD VSS sg13g2_decap_8
X_1621_ _1639_/A _1621_/B _1621_/Y VDD VSS sg13g2_nor2_1
XFILLER_99_625 VDD VSS sg13g2_decap_8
X_1552_ _1551_/Y VDD _1552_/Y VSS _1573_/A1 _2206_/Q sg13g2_o21ai_1
XFILLER_28_1029 VDD VSS sg13g2_decap_8
X_1483_ VDD _2260_/D _1483_/A VSS sg13g2_inv_1
XFILLER_4_581 VDD VSS sg13g2_decap_8
XFILLER_101_608 VDD VSS sg13g2_decap_8
XFILLER_86_308 VDD VSS sg13g2_fill_1
XFILLER_97_91 VDD VSS sg13g2_decap_8
XFILLER_67_511 VDD VSS sg13g2_decap_8
XFILLER_39_224 VDD VSS sg13g2_decap_8
XFILLER_95_875 VDD VSS sg13g2_decap_8
XFILLER_55_706 VDD VSS sg13g2_decap_8
X_2104_ _2106_/B _2104_/B _2094_/B VDD VSS sg13g2_nand2b_1
XFILLER_36_931 VDD VSS sg13g2_decap_8
XFILLER_67_588 VDD VSS sg13g2_decap_8
XFILLER_54_227 VDD VSS sg13g2_fill_2
X_2035_ _2030_/Y VDD _2325_/D VSS _2031_/Y _2034_/Y sg13g2_o21ai_1
XFILLER_82_569 VDD VSS sg13g2_decap_8
XFILLER_35_441 VDD VSS sg13g2_decap_8
XFILLER_63_772 VDD VSS sg13g2_decap_8
XFILLER_74_1038 VDD VSS sg13g2_decap_8
XFILLER_51_989 VDD VSS sg13g2_decap_8
XFILLER_23_658 VDD VSS sg13g2_decap_8
XFILLER_10_308 VDD VSS sg13g2_decap_8
XFILLER_50_444 VDD VSS sg13g2_decap_8
XFILLER_22_168 VDD VSS sg13g2_decap_8
XFILLER_108_207 VDD VSS sg13g2_decap_8
XFILLER_108_229 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[7\].out_data_pad out_data_PADs[7] bondpad_70x70
XFILLER_11_1022 VDD VSS sg13g2_decap_8
XFILLER_105_903 VDD VSS sg13g2_decap_8
X_1819_ _1821_/B _1819_/B _1949_/A VDD VSS sg13g2_nand2b_1
Xhold320 _2179_/Q VDD VSS hold320/X sg13g2_dlygate4sd3_1
Xhold353 _2202_/Q VDD VSS hold353/X sg13g2_dlygate4sd3_1
Xhold342 _1488_/Y VDD VSS _2264_/D sg13g2_dlygate4sd3_1
Xhold331 _2106_/Y VDD VSS _2353_/D sg13g2_dlygate4sd3_1
XFILLER_2_518 VDD VSS sg13g2_decap_8
Xhold375 _2169_/Q VDD VSS hold375/X sg13g2_dlygate4sd3_1
Xhold386 _1308_/Y VDD VSS _1309_/A sg13g2_dlygate4sd3_1
Xhold364 _2182_/Q VDD VSS hold364/X sg13g2_dlygate4sd3_1
XFILLER_77_28 VDD VSS sg13g2_decap_8
XFILLER_89_168 VDD VSS sg13g2_decap_8
XFILLER_89_179 VDD VSS sg13g2_decap_8
XFILLER_77_308 VDD VSS sg13g2_decap_8
Xhold397 _1446_/Y VDD VSS _2243_/D sg13g2_dlygate4sd3_1
XFILLER_98_691 VDD VSS sg13g2_fill_2
XFILLER_58_511 VDD VSS sg13g2_decap_8
XFILLER_100_630 VDD VSS sg13g2_decap_8
XFILLER_112_490 VDD VSS sg13g2_decap_8
XFILLER_85_341 VDD VSS sg13g2_decap_8
XFILLER_58_577 VDD VSS sg13g2_fill_2
XFILLER_100_696 VDD VSS sg13g2_decap_8
XFILLER_39_780 VDD VSS sg13g2_decap_8
XFILLER_93_49 VDD VSS sg13g2_decap_8
XFILLER_27_931 VDD VSS sg13g2_decap_8
XFILLER_26_21 VDD VSS sg13g2_decap_8
XFILLER_54_772 VDD VSS sg13g2_fill_1
XFILLER_26_441 VDD VSS sg13g2_decap_8
XFILLER_81_580 VDD VSS sg13g2_decap_8
XFILLER_42_945 VDD VSS sg13g2_decap_8
XFILLER_26_98 VDD VSS sg13g2_decap_8
XFILLER_14_658 VDD VSS sg13g2_decap_8
XFILLER_41_444 VDD VSS sg13g2_decap_8
XFILLER_13_168 VDD VSS sg13g2_decap_8
XFILLER_42_42 VDD VSS sg13g2_decap_8
XFILLER_5_301 VDD VSS sg13g2_decap_8
XFILLER_10_875 VDD VSS sg13g2_decap_8
XFILLER_108_752 VDD VSS sg13g2_decap_8
X_2327__201 VDD VSS _2327_/RESET_B sg13g2_tiehi
X_2366__261 VDD VSS _2366_/RESET_B sg13g2_tiehi
XFILLER_6_868 VDD VSS sg13g2_decap_8
XFILLER_107_273 VDD VSS sg13g2_decap_4
XFILLER_5_378 VDD VSS sg13g2_decap_8
XFILLER_69_809 VDD VSS sg13g2_decap_8
XFILLER_111_917 VDD VSS sg13g2_decap_8
XFILLER_95_105 VDD VSS sg13g2_decap_8
XFILLER_68_319 VDD VSS sg13g2_decap_8
XFILLER_3_14 VDD VSS sg13g2_decap_8
XFILLER_49_500 VDD VSS sg13g2_decap_8
XFILLER_110_438 VDD VSS sg13g2_decap_8
XFILLER_1_595 VDD VSS sg13g2_decap_8
XFILLER_49_544 VDD VSS sg13g2_decap_8
XFILLER_97_1005 VDD VSS sg13g2_decap_4
XFILLER_92_812 VDD VSS sg13g2_decap_8
XFILLER_37_728 VDD VSS sg13g2_decap_8
XFILLER_64_536 VDD VSS sg13g2_decap_8
XFILLER_18_931 VDD VSS sg13g2_decap_8
XFILLER_36_238 VDD VSS sg13g2_decap_8
XFILLER_91_355 VDD VSS sg13g2_decap_8
XFILLER_45_772 VDD VSS sg13g2_decap_4
XFILLER_45_783 VDD VSS sg13g2_decap_8
XFILLER_17_441 VDD VSS sg13g2_decap_8
XFILLER_72_591 VDD VSS sg13g2_decap_8
XFILLER_33_945 VDD VSS sg13g2_decap_8
XFILLER_32_455 VDD VSS sg13g2_decap_8
XFILLER_73_1060 VDD VSS sg13g2_fill_1
XFILLER_34_1022 VDD VSS sg13g2_decap_8
XFILLER_9_651 VDD VSS sg13g2_decap_8
XFILLER_8_161 VDD VSS sg13g2_decap_8
XFILLER_99_400 VDD VSS sg13g2_decap_4
X_1604_ _1639_/A _1604_/B _1604_/Y VDD VSS sg13g2_nor2_1
X_1535_ _1556_/S0 _2236_/Q _2228_/Q _2220_/Q _2212_/Q _1589_/B _1536_/A VDD VSS sg13g2_mux4_1
XFILLER_99_455 VDD VSS sg13g2_decap_8
XFILLER_101_416 VDD VSS sg13g2_decap_8
X_1466_ _1367_/A VDD _1466_/Y VSS _1364_/A _1481_/A2 sg13g2_o21ai_1
XFILLER_83_801 VDD VSS sg13g2_decap_8
X_1397_ _1398_/A _1392_/Y hold513/X _1392_/B _1373_/A VDD VSS sg13g2_a22oi_1
XFILLER_95_672 VDD VSS sg13g2_decap_8
XFILLER_68_897 VDD VSS sg13g2_decap_8
XFILLER_28_728 VDD VSS sg13g2_decap_8
XFILLER_83_845 VDD VSS sg13g2_fill_1
XFILLER_43_709 VDD VSS sg13g2_decap_8
XFILLER_55_536 VDD VSS sg13g2_decap_4
XFILLER_27_238 VDD VSS sg13g2_decap_8
X_2018_ _2017_/Y VDD _2322_/D VSS _2025_/A _2015_/Y sg13g2_o21ai_1
XFILLER_83_878 VDD VSS sg13g2_decap_8
XFILLER_42_219 VDD VSS sg13g2_decap_8
XFILLER_24_945 VDD VSS sg13g2_decap_8
XFILLER_63_580 VDD VSS sg13g2_fill_1
XFILLER_23_455 VDD VSS sg13g2_decap_8
XFILLER_51_786 VDD VSS sg13g2_decap_8
XFILLER_10_105 VDD VSS sg13g2_decap_8
XFILLER_50_252 VDD VSS sg13g2_decap_8
X_2166__208 VDD VSS _2166_/RESET_B sg13g2_tiehi
XFILLER_12_56 VDD VSS sg13g2_decap_8
XFILLER_105_700 VDD VSS sg13g2_decap_8
XFILLER_3_805 VDD VSS sg13g2_decap_8
XFILLER_88_49 VDD VSS sg13g2_decap_8
XFILLER_2_315 VDD VSS sg13g2_decap_8
XFILLER_105_777 VDD VSS sg13g2_decap_8
XFILLER_78_628 VDD VSS sg13g2_decap_8
XFILLER_104_287 VDD VSS sg13g2_fill_1
XFILLER_77_105 VDD VSS sg13g2_decap_8
XFILLER_58_330 VDD VSS sg13g2_decap_8
XFILLER_86_672 VDD VSS sg13g2_decap_8
XFILLER_100_471 VDD VSS sg13g2_decap_4
XFILLER_58_385 VDD VSS sg13g2_decap_8
XFILLER_19_728 VDD VSS sg13g2_decap_8
XFILLER_37_42 VDD VSS sg13g2_decap_8
XFILLER_46_503 VDD VSS sg13g2_decap_8
XFILLER_74_856 VDD VSS sg13g2_decap_8
XFILLER_85_171 VDD VSS sg13g2_decap_8
XFILLER_73_344 VDD VSS sg13g2_decap_8
XFILLER_18_238 VDD VSS sg13g2_decap_8
XFILLER_57_1000 VDD VSS sg13g2_decap_4
XFILLER_96_1060 VDD VSS sg13g2_fill_1
XFILLER_15_945 VDD VSS sg13g2_decap_8
XFILLER_42_742 VDD VSS sg13g2_decap_8
XFILLER_14_455 VDD VSS sg13g2_decap_8
XFILLER_41_241 VDD VSS sg13g2_decap_8
XFILLER_41_274 VDD VSS sg13g2_decap_8
XFILLER_30_959 VDD VSS sg13g2_decap_8
XFILLER_10_672 VDD VSS sg13g2_decap_8
XFILLER_6_665 VDD VSS sg13g2_decap_8
XFILLER_5_175 VDD VSS sg13g2_decap_8
XFILLER_45_7 VDD VSS sg13g2_decap_8
XFILLER_111_714 VDD VSS sg13g2_decap_8
X_1320_ _1320_/Y _1322_/B1 hold306/X _1322_/A2 _2323_/Q VDD VSS sg13g2_a22oi_1
XFILLER_97_948 VDD VSS sg13g2_fill_1
XFILLER_97_937 VDD VSS sg13g2_decap_8
XFILLER_69_628 VDD VSS sg13g2_decap_8
XFILLER_110_224 VDD VSS sg13g2_decap_8
XFILLER_2_882 VDD VSS sg13g2_decap_8
XFILLER_96_469 VDD VSS sg13g2_decap_4
XFILLER_1_392 VDD VSS sg13g2_decap_8
X_1251_ VSS VDD _2092_/A _2093_/B _1251_/Y _2101_/A sg13g2_a21oi_1
XFILLER_49_330 VDD VSS sg13g2_decap_8
XFILLER_83_119 VDD VSS sg13g2_decap_8
XFILLER_65_834 VDD VSS sg13g2_decap_8
XFILLER_64_300 VDD VSS sg13g2_decap_8
XFILLER_37_525 VDD VSS sg13g2_decap_8
X_2305__91 VDD VSS _2305__91/L_HI sg13g2_tiehi
XFILLER_76_182 VDD VSS sg13g2_decap_8
XFILLER_94_70 VDD VSS sg13g2_decap_8
XFILLER_65_845 VDD VSS sg13g2_fill_2
XFILLER_92_675 VDD VSS sg13g2_decap_8
XFILLER_64_388 VDD VSS sg13g2_decap_8
XFILLER_33_742 VDD VSS sg13g2_decap_8
XFILLER_71_1019 VDD VSS sg13g2_decap_8
XFILLER_32_252 VDD VSS sg13g2_decap_8
XFILLER_21_959 VDD VSS sg13g2_decap_8
XFILLER_71_0 VDD VSS sg13g2_decap_8
XFILLER_20_469 VDD VSS sg13g2_decap_8
XFILLER_99_263 VDD VSS sg13g2_decap_8
XFILLER_0_819 VDD VSS sg13g2_decap_8
XFILLER_102_714 VDD VSS sg13g2_fill_1
XFILLER_101_213 VDD VSS sg13g2_decap_8
X_1518_ _1518_/B _1518_/C _2273_/Q _1518_/Y VDD VSS _1518_/D sg13g2_nand4_1
XFILLER_75_609 VDD VSS sg13g2_decap_8
XFILLER_87_458 VDD VSS sg13g2_decap_4
X_1449_ _1449_/A _1463_/B _1449_/Y VDD VSS sg13g2_nor2_1
XFILLER_96_992 VDD VSS sg13g2_decap_8
XFILLER_74_119 VDD VSS sg13g2_decap_8
XFILLER_56_812 VDD VSS sg13g2_decap_4
XFILLER_67_160 VDD VSS sg13g2_decap_8
XFILLER_68_694 VDD VSS sg13g2_decap_8
XFILLER_55_322 VDD VSS sg13g2_decap_8
XFILLER_28_525 VDD VSS sg13g2_decap_8
XFILLER_71_826 VDD VSS sg13g2_decap_8
XFILLER_56_878 VDD VSS sg13g2_decap_8
XFILLER_55_355 VDD VSS sg13g2_fill_2
XFILLER_55_377 VDD VSS sg13g2_fill_2
XFILLER_82_163 VDD VSS sg13g2_decap_8
XFILLER_55_399 VDD VSS sg13g2_decap_8
XFILLER_43_539 VDD VSS sg13g2_fill_2
XFILLER_43_528 VDD VSS sg13g2_decap_8
XFILLER_70_358 VDD VSS sg13g2_decap_8
XFILLER_90_28 VDD VSS sg13g2_decap_8
XFILLER_24_742 VDD VSS sg13g2_decap_8
XFILLER_51_572 VDD VSS sg13g2_decap_8
XFILLER_23_252 VDD VSS sg13g2_decap_8
XFILLER_12_959 VDD VSS sg13g2_decap_8
XFILLER_17_1050 VDD VSS sg13g2_decap_8
XFILLER_104_1020 VDD VSS sg13g2_decap_8
XFILLER_11_469 VDD VSS sg13g2_decap_8
XFILLER_23_77 VDD VSS sg13g2_decap_8
XFILLER_87_1004 VDD VSS sg13g2_decap_8
XFILLER_109_324 VDD VSS sg13g2_fill_1
XFILLER_3_602 VDD VSS sg13g2_decap_8
Xout_ready_pad IOVDD IOVSS _1259_/C out_ready_PAD VDD VSS sg13g2_IOPadIn
XFILLER_2_112 VDD VSS sg13g2_decap_8
XFILLER_78_403 VDD VSS sg13g2_decap_8
XFILLER_3_679 VDD VSS sg13g2_decap_8
XFILLER_105_574 VDD VSS sg13g2_decap_8
XFILLER_2_189 VDD VSS sg13g2_decap_8
XFILLER_93_428 VDD VSS sg13g2_decap_8
XFILLER_24_1043 VDD VSS sg13g2_decap_8
XFILLER_48_63 VDD VSS sg13g2_decap_8
XFILLER_65_108 VDD VSS sg13g2_decap_4
XFILLER_47_845 VDD VSS sg13g2_fill_1
XFILLER_19_525 VDD VSS sg13g2_decap_8
XFILLER_46_333 VDD VSS sg13g2_decap_8
XFILLER_111_1057 VDD VSS sg13g2_decap_4
XFILLER_74_653 VDD VSS sg13g2_decap_8
XFILLER_73_130 VDD VSS sg13g2_fill_1
XFILLER_73_185 VDD VSS sg13g2_decap_4
XFILLER_104_91 VDD VSS sg13g2_decap_8
XFILLER_34_539 VDD VSS sg13g2_decap_8
XFILLER_61_347 VDD VSS sg13g2_decap_8
XFILLER_15_742 VDD VSS sg13g2_decap_8
XFILLER_70_892 VDD VSS sg13g2_decap_8
XFILLER_14_252 VDD VSS sg13g2_decap_8
XFILLER_9_35 VDD VSS sg13g2_decap_8
XFILLER_30_756 VDD VSS sg13g2_decap_8
XFILLER_31_1036 VDD VSS sg13g2_decap_8
XFILLER_7_952 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_6_462 VDD VSS sg13g2_decap_8
XFILLER_89_70 VDD VSS sg13g2_decap_8
XFILLER_111_511 VDD VSS sg13g2_decap_8
XFILLER_69_414 VDD VSS sg13g2_fill_2
XFILLER_9_1015 VDD VSS sg13g2_decap_8
X_2352_ _2352__89/L_HI VSS VDD _2352_/D _2352_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_97_778 VDD VSS sg13g2_decap_8
XFILLER_85_907 VDD VSS sg13g2_decap_8
X_1303_ VDD _2181_/D _1303_/A VSS sg13g2_inv_1
X_2283_ _2283_/RESET_B VSS VDD _2283_/D _2283_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_85_929 VDD VSS sg13g2_decap_8
XFILLER_111_588 VDD VSS sg13g2_decap_8
XFILLER_96_266 VDD VSS sg13g2_decap_8
X_1234_ _1235_/A _1234_/B _1492_/B VDD VSS sg13g2_nor2_1
XFILLER_93_951 VDD VSS sg13g2_decap_8
XFILLER_84_439 VDD VSS sg13g2_fill_1
XFILLER_38_856 VDD VSS sg13g2_decap_8
XFILLER_37_322 VDD VSS sg13g2_decap_8
XFILLER_49_182 VDD VSS sg13g2_decap_8
XFILLER_65_675 VDD VSS sg13g2_decap_8
XFILLER_80_623 VDD VSS sg13g2_decap_8
XFILLER_53_859 VDD VSS sg13g2_decap_8
XFILLER_25_539 VDD VSS sg13g2_decap_8
XFILLER_37_399 VDD VSS sg13g2_decap_8
XFILLER_80_678 VDD VSS sg13g2_decap_8
XFILLER_100_49 VDD VSS sg13g2_decap_8
XFILLER_21_756 VDD VSS sg13g2_decap_8
XFILLER_60_391 VDD VSS sg13g2_decap_8
XFILLER_20_266 VDD VSS sg13g2_decap_8
X_1998_ _1999_/A _2021_/S _1998_/X VDD VSS sg13g2_and2_1
XFILLER_109_14 VDD VSS sg13g2_decap_8
XFILLER_107_828 VDD VSS sg13g2_decap_8
XFILLER_106_305 VDD VSS sg13g2_decap_8
XFILLER_0_616 VDD VSS sg13g2_decap_8
XFILLER_76_918 VDD VSS sg13g2_fill_1
XFILLER_88_767 VDD VSS sg13g2_decap_8
XFILLER_76_907 VDD VSS sg13g2_decap_8
XFILLER_87_222 VDD VSS sg13g2_decap_8
XFILLER_87_233 VDD VSS sg13g2_decap_4
XFILLER_102_588 VDD VSS sg13g2_decap_8
XFILLER_87_255 VDD VSS sg13g2_decap_8
XFILLER_85_28 VDD VSS sg13g2_decap_8
XFILLER_29_812 VDD VSS sg13g2_decap_8
XFILLER_68_480 VDD VSS sg13g2_decap_8
XFILLER_28_322 VDD VSS sg13g2_decap_8
XFILLER_84_973 VDD VSS sg13g2_decap_8
XFILLER_44_804 VDD VSS sg13g2_decap_8
XFILLER_29_889 VDD VSS sg13g2_decap_8
XFILLER_18_77 VDD VSS sg13g2_decap_8
XFILLER_71_612 VDD VSS sg13g2_decap_8
XFILLER_83_494 VDD VSS sg13g2_fill_1
XFILLER_16_539 VDD VSS sg13g2_decap_8
XFILLER_28_399 VDD VSS sg13g2_decap_8
XFILLER_70_133 VDD VSS sg13g2_decap_8
XFILLER_55_196 VDD VSS sg13g2_decap_8
XFILLER_34_21 VDD VSS sg13g2_decap_8
XFILLER_43_336 VDD VSS sg13g2_decap_8
XFILLER_93_1052 VDD VSS sg13g2_decap_8
XFILLER_52_870 VDD VSS sg13g2_decap_4
XFILLER_54_1036 VDD VSS sg13g2_decap_8
XFILLER_12_756 VDD VSS sg13g2_decap_8
XFILLER_34_98 VDD VSS sg13g2_decap_8
XFILLER_11_266 VDD VSS sg13g2_decap_8
XFILLER_8_749 VDD VSS sg13g2_decap_8
XFILLER_109_154 VDD VSS sg13g2_decap_8
XFILLER_7_259 VDD VSS sg13g2_decap_8
XFILLER_50_86 VDD VSS sg13g2_fill_2
XFILLER_4_966 VDD VSS sg13g2_decap_8
XFILLER_112_308 VDD VSS sg13g2_decap_8
XFILLER_3_476 VDD VSS sg13g2_decap_8
XFILLER_1_0 VDD VSS sg13g2_decap_8
XFILLER_105_393 VDD VSS sg13g2_decap_8
XFILLER_79_778 VDD VSS sg13g2_decap_8
XFILLER_66_417 VDD VSS sg13g2_fill_2
XFILLER_66_428 VDD VSS sg13g2_decap_8
XFILLER_66_406 VDD VSS sg13g2_decap_8
XFILLER_38_119 VDD VSS sg13g2_decap_8
XFILLER_19_322 VDD VSS sg13g2_decap_8
X_2294__133 VDD VSS _2294_/RESET_B sg13g2_tiehi
XFILLER_74_461 VDD VSS sg13g2_decap_8
XFILLER_35_826 VDD VSS sg13g2_decap_8
XFILLER_19_399 VDD VSS sg13g2_decap_8
XFILLER_46_185 VDD VSS sg13g2_decap_8
XFILLER_34_336 VDD VSS sg13g2_decap_8
XFILLER_90_987 VDD VSS sg13g2_decap_8
X_2335__163 VDD VSS _2335_/RESET_B sg13g2_tiehi
XFILLER_43_870 VDD VSS sg13g2_decap_8
X_1921_ _1921_/Y _1921_/A _1921_/B VDD VSS sg13g2_xnor2_1
XFILLER_61_199 VDD VSS sg13g2_decap_8
XFILLER_42_391 VDD VSS sg13g2_decap_8
XFILLER_30_553 VDD VSS sg13g2_decap_8
X_1852_ _1852_/B _1852_/C _1852_/A _1866_/A VDD VSS sg13g2_nand3_1
X_1783_ _1929_/B _2212_/Q _2220_/Q VDD VSS sg13g2_xnor2_1
Xfanout9 _2061_/S _2079_/S VDD VSS sg13g2_buf_1
XFILLER_69_211 VDD VSS sg13g2_decap_8
XFILLER_97_542 VDD VSS sg13g2_decap_8
XFILLER_34_0 VDD VSS sg13g2_decap_8
XFILLER_112_875 VDD VSS sg13g2_decap_8
XFILLER_85_715 VDD VSS sg13g2_fill_2
XFILLER_58_929 VDD VSS sg13g2_decap_8
X_2335_ _2335_/RESET_B VSS VDD _2335_/D _2335_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_111_385 VDD VSS sg13g2_decap_8
XFILLER_84_214 VDD VSS sg13g2_decap_8
XFILLER_69_288 VDD VSS sg13g2_decap_8
XFILLER_57_439 VDD VSS sg13g2_decap_8
X_2266_ _2266_/RESET_B VSS VDD _2266_/D _2266_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_29_119 VDD VSS sg13g2_decap_8
X_2197_ _2197_/RESET_B VSS VDD _2197_/D _2197_/Q _2345_/CLK sg13g2_dfrbpq_1
X_1217_ VDD _1726_/A _2234_/Q VSS sg13g2_inv_1
XFILLER_38_653 VDD VSS sg13g2_decap_8
XFILLER_81_932 VDD VSS sg13g2_decap_8
XFILLER_77_1014 VDD VSS sg13g2_decap_8
XFILLER_66_984 VDD VSS sg13g2_fill_1
XFILLER_53_623 VDD VSS sg13g2_decap_8
XFILLER_26_826 VDD VSS sg13g2_decap_8
XFILLER_1_91 VDD VSS sg13g2_decap_8
XFILLER_52_100 VDD VSS sg13g2_fill_2
Xout_data_pads\[4\].out_data_pad _2370_/Q IOVDD IOVSS out_data_PADs[4] VDD VSS sg13g2_IOPadOut30mA
XFILLER_92_291 VDD VSS sg13g2_decap_8
XFILLER_65_494 VDD VSS sg13g2_decap_8
XFILLER_25_336 VDD VSS sg13g2_decap_8
XFILLER_37_196 VDD VSS sg13g2_decap_8
XFILLER_80_453 VDD VSS sg13g2_decap_8
XFILLER_41_818 VDD VSS sg13g2_decap_8
XFILLER_40_328 VDD VSS sg13g2_decap_8
XFILLER_52_188 VDD VSS sg13g2_decap_8
XFILLER_21_553 VDD VSS sg13g2_decap_8
XFILLER_101_1023 VDD VSS sg13g2_decap_8
XFILLER_101_1034 VDD VSS sg13g2_decap_8
XFILLER_107_625 VDD VSS sg13g2_decap_8
XFILLER_112_7 VDD VSS sg13g2_decap_8
XFILLER_20_56 VDD VSS sg13g2_decap_8
XFILLER_1_903 VDD VSS sg13g2_decap_8
XFILLER_106_168 VDD VSS sg13g2_decap_8
XFILLER_0_413 VDD VSS sg13g2_decap_8
XFILLER_96_49 VDD VSS sg13g2_decap_8
X_2360__278 VDD VSS _2360_/RESET_B sg13g2_tiehi
XFILLER_103_886 VDD VSS sg13g2_fill_1
XFILLER_88_575 VDD VSS sg13g2_decap_8
XFILLER_49_918 VDD VSS sg13g2_fill_2
XFILLER_29_21 VDD VSS sg13g2_decap_8
XFILLER_76_748 VDD VSS sg13g2_decap_8
XFILLER_102_396 VDD VSS sg13g2_decap_8
XFILLER_75_236 VDD VSS sg13g2_decap_8
XFILLER_29_98 VDD VSS sg13g2_decap_8
XFILLER_84_792 VDD VSS sg13g2_fill_1
XFILLER_84_781 VDD VSS sg13g2_decap_8
XFILLER_21_1057 VDD VSS sg13g2_decap_4
XFILLER_29_686 VDD VSS sg13g2_decap_8
XFILLER_56_483 VDD VSS sg13g2_decap_8
XFILLER_56_461 VDD VSS sg13g2_decap_8
XFILLER_17_826 VDD VSS sg13g2_decap_8
XFILLER_72_976 VDD VSS sg13g2_decap_8
XFILLER_44_634 VDD VSS sg13g2_decap_4
XFILLER_16_336 VDD VSS sg13g2_decap_8
XFILLER_43_133 VDD VSS sg13g2_decap_8
XFILLER_45_42 VDD VSS sg13g2_decap_8
XFILLER_28_196 VDD VSS sg13g2_decap_8
XFILLER_71_453 VDD VSS sg13g2_decap_8
XFILLER_101_70 VDD VSS sg13g2_decap_8
XFILLER_40_851 VDD VSS sg13g2_decap_8
XFILLER_12_553 VDD VSS sg13g2_decap_8
XFILLER_8_546 VDD VSS sg13g2_decap_8
XFILLER_61_63 VDD VSS sg13g2_decap_8
XFILLER_6_14 VDD VSS sg13g2_decap_8
XFILLER_99_829 VDD VSS sg13g2_decap_8
XFILLER_98_339 VDD VSS sg13g2_decap_8
XFILLER_112_105 VDD VSS sg13g2_decap_8
XFILLER_4_763 VDD VSS sg13g2_decap_8
XFILLER_3_273 VDD VSS sg13g2_decap_8
X_2120_ _2120_/A _2120_/B _2120_/Y VDD VSS sg13g2_nor2_1
XFILLER_67_748 VDD VSS sg13g2_decap_4
XFILLER_0_980 VDD VSS sg13g2_decap_8
XFILLER_6_1029 VDD VSS sg13g2_decap_8
XFILLER_94_556 VDD VSS sg13g2_decap_8
XFILLER_94_567 VDD VSS sg13g2_fill_1
X_2051_ _2049_/X _2050_/X _2079_/S _2077_/A VDD VSS sg13g2_mux2_1
XFILLER_86_93 VDD VSS sg13g2_fill_1
XFILLER_48_951 VDD VSS sg13g2_fill_1
XFILLER_66_258 VDD VSS sg13g2_fill_2
XFILLER_81_217 VDD VSS sg13g2_decap_4
XFILLER_48_995 VDD VSS sg13g2_decap_8
XFILLER_35_623 VDD VSS sg13g2_decap_8
XFILLER_62_442 VDD VSS sg13g2_decap_8
XFILLER_19_196 VDD VSS sg13g2_decap_8
XFILLER_34_133 VDD VSS sg13g2_decap_8
XFILLER_90_773 VDD VSS sg13g2_decap_8
XFILLER_50_604 VDD VSS sg13g2_decap_8
X_1904_ _1905_/A _1905_/B _1920_/B VDD VSS sg13g2_nor2_1
XFILLER_31_840 VDD VSS sg13g2_decap_8
XFILLER_30_350 VDD VSS sg13g2_decap_8
X_1835_ _2205_/Q _2246_/Q _1905_/A VDD VSS sg13g2_xor2_1
X_1766_ _1899_/A _1770_/A _1766_/B VDD VSS sg13g2_nand2_1
Xhold502 _1626_/Y VDD VSS _2294_/D sg13g2_dlygate4sd3_1
Xhold535 _2370_/Q VDD VSS hold535/X sg13g2_dlygate4sd3_1
Xhold513 _2221_/Q VDD VSS hold513/X sg13g2_dlygate4sd3_1
Xhold524 _1610_/Y VDD VSS _2291_/D sg13g2_dlygate4sd3_1
X_1697_ _1703_/A _2315_/Q _1697_/B VDD VSS sg13g2_xnor2_1
XFILLER_89_328 VDD VSS sg13g2_decap_8
XFILLER_103_105 VDD VSS sg13g2_decap_8
Xhold568 _2122_/Y VDD VSS _2367_/D sg13g2_dlygate4sd3_1
Xhold546 _1518_/Y VDD VSS hold546/X sg13g2_dlygate4sd3_1
Xhold557 _2364_/Q VDD VSS _1252_/B sg13g2_dlygate4sd3_1
XFILLER_112_672 VDD VSS sg13g2_decap_8
XFILLER_98_884 VDD VSS sg13g2_decap_8
XFILLER_97_350 VDD VSS sg13g2_fill_2
X_2318_ _2318_/RESET_B VSS VDD _2318_/D _2318_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_111_182 VDD VSS sg13g2_decap_8
XFILLER_97_372 VDD VSS sg13g2_decap_8
XFILLER_73_707 VDD VSS sg13g2_decap_8
XFILLER_39_962 VDD VSS sg13g2_decap_8
XFILLER_57_269 VDD VSS sg13g2_decap_8
XFILLER_45_409 VDD VSS sg13g2_fill_1
XFILLER_85_589 VDD VSS sg13g2_decap_4
XFILLER_72_228 VDD VSS sg13g2_decap_8
XFILLER_26_623 VDD VSS sg13g2_decap_8
X_2249_ _2249_/RESET_B VSS VDD _2249_/D _2249_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_72_239 VDD VSS sg13g2_fill_1
XFILLER_53_442 VDD VSS sg13g2_decap_8
XFILLER_25_133 VDD VSS sg13g2_decap_8
XFILLER_54_976 VDD VSS sg13g2_decap_8
XFILLER_41_615 VDD VSS sg13g2_decap_8
XFILLER_90_1022 VDD VSS sg13g2_decap_8
XFILLER_80_283 VDD VSS sg13g2_decap_8
XFILLER_15_56 VDD VSS sg13g2_decap_8
XFILLER_22_840 VDD VSS sg13g2_decap_8
XFILLER_40_147 VDD VSS sg13g2_decap_8
XFILLER_51_1017 VDD VSS sg13g2_decap_8
XFILLER_21_350 VDD VSS sg13g2_decap_8
XFILLER_108_934 VDD VSS sg13g2_decap_8
XFILLER_31_77 VDD VSS sg13g2_decap_8
XFILLER_107_444 VDD VSS sg13g2_decap_8
XFILLER_1_700 VDD VSS sg13g2_decap_8
XFILLER_0_210 VDD VSS sg13g2_decap_8
XFILLER_89_873 VDD VSS sg13g2_decap_8
XFILLER_49_704 VDD VSS sg13g2_decap_8
XFILLER_1_777 VDD VSS sg13g2_decap_8
XFILLER_103_683 VDD VSS sg13g2_fill_1
XFILLER_103_672 VDD VSS sg13g2_decap_8
XFILLER_88_394 VDD VSS sg13g2_decap_8
XFILLER_76_512 VDD VSS sg13g2_decap_8
XFILLER_0_287 VDD VSS sg13g2_decap_8
XFILLER_102_182 VDD VSS sg13g2_fill_2
XFILLER_64_718 VDD VSS sg13g2_decap_8
XFILLER_76_589 VDD VSS sg13g2_decap_8
XFILLER_45_954 VDD VSS sg13g2_decap_8
XFILLER_63_239 VDD VSS sg13g2_decap_4
XFILLER_56_291 VDD VSS sg13g2_decap_8
XFILLER_17_623 VDD VSS sg13g2_decap_8
XFILLER_29_483 VDD VSS sg13g2_decap_8
XFILLER_72_773 VDD VSS sg13g2_decap_8
XFILLER_16_133 VDD VSS sg13g2_decap_8
XFILLER_44_453 VDD VSS sg13g2_decap_8
XFILLER_108_1018 VDD VSS sg13g2_decap_8
XFILLER_112_91 VDD VSS sg13g2_decap_8
XFILLER_60_935 VDD VSS sg13g2_decap_8
XFILLER_32_637 VDD VSS sg13g2_decap_8
XFILLER_13_840 VDD VSS sg13g2_decap_8
XFILLER_31_147 VDD VSS sg13g2_decap_8
XFILLER_12_350 VDD VSS sg13g2_decap_8
XFILLER_9_833 VDD VSS sg13g2_decap_8
XFILLER_75_7 VDD VSS sg13g2_decap_8
XFILLER_8_343 VDD VSS sg13g2_decap_8
X_1620_ _1619_/Y VDD _1620_/Y VSS _1634_/A hold551/X sg13g2_o21ai_1
X_1551_ VSS VDD _1573_/A1 _1212_/Y _1551_/Y _1523_/B sg13g2_a21oi_1
XFILLER_67_1046 VDD VSS sg13g2_decap_8
XFILLER_28_1008 VDD VSS sg13g2_decap_8
X_2263__227 VDD VSS _2263_/RESET_B sg13g2_tiehi
XFILLER_4_560 VDD VSS sg13g2_decap_8
XFILLER_99_659 VDD VSS sg13g2_decap_8
X_1482_ _1483_/A _1482_/B1 _2110_/B _1482_/A2 _1485_/A VDD VSS sg13g2_a22oi_1
XFILLER_97_70 VDD VSS sg13g2_decap_8
XFILLER_95_843 VDD VSS sg13g2_decap_4
XFILLER_100_119 VDD VSS sg13g2_decap_8
XFILLER_39_203 VDD VSS sg13g2_decap_8
XFILLER_67_567 VDD VSS sg13g2_decap_8
X_2103_ VDD _2103_/Y _2104_/B VSS sg13g2_inv_1
XFILLER_36_910 VDD VSS sg13g2_decap_8
X_2034_ _2034_/Y _2082_/B _2034_/B VDD VSS sg13g2_nand2_1
XFILLER_82_548 VDD VSS sg13g2_decap_8
XFILLER_35_420 VDD VSS sg13g2_decap_8
XFILLER_74_1017 VDD VSS sg13g2_decap_8
XFILLER_36_987 VDD VSS sg13g2_decap_8
XFILLER_63_751 VDD VSS sg13g2_decap_8
XFILLER_90_570 VDD VSS sg13g2_decap_8
XFILLER_90_581 VDD VSS sg13g2_fill_2
XFILLER_51_946 VDD VSS sg13g2_fill_2
XFILLER_23_637 VDD VSS sg13g2_decap_8
XFILLER_35_497 VDD VSS sg13g2_decap_8
XFILLER_50_423 VDD VSS sg13g2_decap_8
XFILLER_62_294 VDD VSS sg13g2_decap_4
XFILLER_22_147 VDD VSS sg13g2_decap_8
X_1818_ VSS VDD _1809_/A _1809_/B _1949_/B _1819_/B sg13g2_a21oi_1
XFILLER_11_1001 VDD VSS sg13g2_decap_8
Xhold310 _2173_/Q VDD VSS hold310/X sg13g2_dlygate4sd3_1
Xhold343 _2192_/Q VDD VSS hold343/X sg13g2_dlygate4sd3_1
Xhold332 _2178_/Q VDD VSS hold332/X sg13g2_dlygate4sd3_1
X_1749_ _1749_/A _1751_/B _1762_/A VDD VSS sg13g2_nor2b_1
XFILLER_104_403 VDD VSS sg13g2_fill_2
Xhold321 _1298_/Y VDD VSS _1299_/A sg13g2_dlygate4sd3_1
XFILLER_105_959 VDD VSS sg13g2_decap_8
Xhold376 _1278_/Y VDD VSS _1279_/A sg13g2_dlygate4sd3_1
Xhold387 _2183_/Q VDD VSS hold387/X sg13g2_dlygate4sd3_1
Xhold365 _1304_/Y VDD VSS _1305_/A sg13g2_dlygate4sd3_1
Xhold354 _1344_/Y VDD VSS _1345_/A sg13g2_dlygate4sd3_1
XFILLER_104_458 VDD VSS sg13g2_decap_8
XFILLER_89_147 VDD VSS sg13g2_decap_8
Xhold398 _2253_/Q VDD VSS _1200_/A sg13g2_dlygate4sd3_1
XFILLER_98_670 VDD VSS sg13g2_decap_8
XFILLER_86_876 VDD VSS sg13g2_decap_8
XFILLER_85_320 VDD VSS sg13g2_decap_8
XFILLER_100_675 VDD VSS sg13g2_decap_8
XFILLER_93_28 VDD VSS sg13g2_decap_8
XFILLER_27_910 VDD VSS sg13g2_decap_8
XFILLER_45_217 VDD VSS sg13g2_decap_4
XFILLER_85_397 VDD VSS sg13g2_decap_8
XFILLER_26_420 VDD VSS sg13g2_decap_8
XFILLER_38_280 VDD VSS sg13g2_decap_8
XFILLER_27_987 VDD VSS sg13g2_decap_8
XFILLER_54_751 VDD VSS sg13g2_decap_8
XFILLER_42_924 VDD VSS sg13g2_decap_8
XFILLER_14_637 VDD VSS sg13g2_decap_8
XFILLER_26_77 VDD VSS sg13g2_decap_8
XFILLER_26_497 VDD VSS sg13g2_decap_8
XFILLER_41_423 VDD VSS sg13g2_decap_8
XFILLER_13_147 VDD VSS sg13g2_decap_8
XFILLER_41_467 VDD VSS sg13g2_fill_1
XFILLER_42_21 VDD VSS sg13g2_decap_8
XFILLER_10_854 VDD VSS sg13g2_decap_8
XFILLER_42_98 VDD VSS sg13g2_decap_8
XFILLER_108_731 VDD VSS sg13g2_decap_8
XFILLER_6_847 VDD VSS sg13g2_decap_8
XFILLER_107_252 VDD VSS sg13g2_decap_8
XFILLER_101_0 VDD VSS sg13g2_decap_8
XFILLER_5_357 VDD VSS sg13g2_decap_8
XFILLER_104_992 VDD VSS sg13g2_decap_8
XFILLER_89_692 VDD VSS sg13g2_decap_8
XFILLER_110_417 VDD VSS sg13g2_decap_8
XFILLER_107_91 VDD VSS sg13g2_decap_8
XFILLER_1_574 VDD VSS sg13g2_decap_8
XFILLER_76_331 VDD VSS sg13g2_decap_8
XFILLER_37_707 VDD VSS sg13g2_decap_8
XFILLER_67_84 VDD VSS sg13g2_decap_8
XFILLER_77_898 VDD VSS sg13g2_decap_8
XFILLER_64_515 VDD VSS sg13g2_decap_8
XFILLER_18_910 VDD VSS sg13g2_decap_8
XFILLER_36_217 VDD VSS sg13g2_decap_8
XFILLER_92_868 VDD VSS sg13g2_decap_4
XFILLER_91_334 VDD VSS sg13g2_decap_8
XFILLER_17_420 VDD VSS sg13g2_decap_8
XFILLER_29_280 VDD VSS sg13g2_decap_8
XFILLER_45_751 VDD VSS sg13g2_decap_8
XFILLER_18_987 VDD VSS sg13g2_decap_8
XFILLER_51_209 VDD VSS sg13g2_decap_8
XFILLER_72_570 VDD VSS sg13g2_decap_8
XFILLER_91_389 VDD VSS sg13g2_decap_8
XFILLER_33_924 VDD VSS sg13g2_decap_8
XFILLER_17_497 VDD VSS sg13g2_decap_8
XFILLER_44_272 VDD VSS sg13g2_decap_8
XFILLER_44_261 VDD VSS sg13g2_fill_1
XFILLER_60_743 VDD VSS sg13g2_fill_1
XFILLER_32_434 VDD VSS sg13g2_decap_8
XFILLER_44_294 VDD VSS sg13g2_decap_8
XFILLER_34_1001 VDD VSS sg13g2_decap_8
XFILLER_9_630 VDD VSS sg13g2_decap_8
XFILLER_8_140 VDD VSS sg13g2_decap_8
X_1603_ _1601_/Y VDD _1603_/Y VSS _1638_/S hold527/X sg13g2_o21ai_1
X_1534_ _1576_/A _1534_/B _2275_/D VDD VSS sg13g2_nor2_1
XIO_FILL_IO_EAST_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_80_1043 VDD VSS sg13g2_decap_8
X_1465_ _1465_/B _1465_/C _2267_/Q _1465_/Y VDD VSS sg13g2_nand3_1
XFILLER_95_651 VDD VSS sg13g2_decap_8
X_1396_ VDD _2220_/D _1396_/A VSS sg13g2_inv_1
XFILLER_68_876 VDD VSS sg13g2_decap_8
XFILLER_28_707 VDD VSS sg13g2_decap_8
XFILLER_110_984 VDD VSS sg13g2_decap_8
XFILLER_94_161 VDD VSS sg13g2_fill_1
XFILLER_41_1049 VDD VSS sg13g2_decap_8
XFILLER_67_364 VDD VSS sg13g2_decap_4
XFILLER_55_515 VDD VSS sg13g2_decap_8
XFILLER_27_217 VDD VSS sg13g2_decap_8
XFILLER_83_857 VDD VSS sg13g2_decap_8
XFILLER_103_49 VDD VSS sg13g2_decap_8
X_2017_ _2017_/Y _2074_/A _2017_/B VDD VSS sg13g2_nand2_1
XFILLER_24_924 VDD VSS sg13g2_decap_8
XFILLER_51_710 VDD VSS sg13g2_decap_8
XFILLER_36_784 VDD VSS sg13g2_decap_8
XFILLER_51_765 VDD VSS sg13g2_decap_8
XFILLER_23_434 VDD VSS sg13g2_decap_8
XFILLER_35_294 VDD VSS sg13g2_decap_8
XFILLER_50_231 VDD VSS sg13g2_decap_8
XFILLER_50_297 VDD VSS sg13g2_decap_8
XFILLER_109_539 VDD VSS sg13g2_decap_8
XFILLER_12_35 VDD VSS sg13g2_decap_8
XFILLER_88_28 VDD VSS sg13g2_decap_8
XFILLER_5_7 VDD VSS sg13g2_decap_8
XFILLER_105_756 VDD VSS sg13g2_decap_8
X_2281__179 VDD VSS _2281_/RESET_B sg13g2_tiehi
XFILLER_104_266 VDD VSS sg13g2_decap_8
XFILLER_59_810 VDD VSS sg13g2_decap_8
XFILLER_101_984 VDD VSS sg13g2_decap_8
XFILLER_101_995 VDD VSS sg13g2_decap_8
XFILLER_85_150 VDD VSS sg13g2_decap_8
XFILLER_19_707 VDD VSS sg13g2_decap_8
XFILLER_37_21 VDD VSS sg13g2_decap_8
XFILLER_74_835 VDD VSS sg13g2_decap_8
XFILLER_18_217 VDD VSS sg13g2_decap_8
XFILLER_46_537 VDD VSS sg13g2_decap_8
XFILLER_2_1043 VDD VSS sg13g2_decap_8
XFILLER_37_98 VDD VSS sg13g2_decap_8
XFILLER_42_721 VDD VSS sg13g2_decap_8
XFILLER_27_784 VDD VSS sg13g2_decap_8
XFILLER_61_529 VDD VSS sg13g2_decap_8
XFILLER_15_924 VDD VSS sg13g2_decap_8
XFILLER_14_434 VDD VSS sg13g2_decap_8
XFILLER_18_1029 VDD VSS sg13g2_decap_8
XFILLER_26_294 VDD VSS sg13g2_decap_8
XFILLER_30_938 VDD VSS sg13g2_decap_8
XFILLER_42_798 VDD VSS sg13g2_decap_8
XFILLER_53_97 VDD VSS sg13g2_decap_8
XFILLER_10_651 VDD VSS sg13g2_decap_8
XFILLER_6_644 VDD VSS sg13g2_decap_8
XFILLER_5_154 VDD VSS sg13g2_decap_8
XFILLER_97_916 VDD VSS sg13g2_decap_8
XFILLER_69_607 VDD VSS sg13g2_decap_8
XFILLER_2_861 VDD VSS sg13g2_decap_8
XFILLER_110_203 VDD VSS sg13g2_decap_8
XFILLER_64_1049 VDD VSS sg13g2_decap_8
XFILLER_1_371 VDD VSS sg13g2_decap_8
XFILLER_38_7 VDD VSS sg13g2_decap_8
XFILLER_68_117 VDD VSS sg13g2_decap_8
XFILLER_96_448 VDD VSS sg13g2_decap_8
X_1250_ _2093_/B _1501_/B _1250_/B VDD VSS sg13g2_nand2_1
XFILLER_76_161 VDD VSS sg13g2_decap_8
XFILLER_65_813 VDD VSS sg13g2_decap_8
XFILLER_37_504 VDD VSS sg13g2_decap_8
XFILLER_92_621 VDD VSS sg13g2_decap_8
XFILLER_77_695 VDD VSS sg13g2_decap_8
XFILLER_92_654 VDD VSS sg13g2_decap_8
XFILLER_64_367 VDD VSS sg13g2_decap_8
XFILLER_91_164 VDD VSS sg13g2_decap_8
XFILLER_45_581 VDD VSS sg13g2_decap_8
XFILLER_33_721 VDD VSS sg13g2_decap_8
XFILLER_18_784 VDD VSS sg13g2_decap_8
XFILLER_17_294 VDD VSS sg13g2_decap_8
XFILLER_32_231 VDD VSS sg13g2_decap_8
XFILLER_21_938 VDD VSS sg13g2_decap_8
XFILLER_60_573 VDD VSS sg13g2_decap_8
XFILLER_33_798 VDD VSS sg13g2_decap_8
XFILLER_20_448 VDD VSS sg13g2_decap_8
XFILLER_64_0 VDD VSS sg13g2_decap_8
XFILLER_99_242 VDD VSS sg13g2_decap_8
XFILLER_87_437 VDD VSS sg13g2_decap_8
X_1517_ VSS VDD _1515_/Y _1516_/X _1517_/Y _1228_/A sg13g2_a21oi_1
XFILLER_59_117 VDD VSS sg13g2_decap_8
XFILLER_99_297 VDD VSS sg13g2_decap_8
X_1448_ _1493_/A _2267_/Q _1583_/A _1448_/X VDD VSS sg13g2_a21o_1
XFILLER_4_91 VDD VSS sg13g2_decap_8
XFILLER_96_971 VDD VSS sg13g2_decap_8
XFILLER_101_269 VDD VSS sg13g2_decap_8
XFILLER_68_673 VDD VSS sg13g2_decap_8
X_2202__136 VDD VSS _2202_/RESET_B sg13g2_tiehi
XFILLER_55_301 VDD VSS sg13g2_decap_8
XFILLER_28_504 VDD VSS sg13g2_decap_8
XFILLER_110_781 VDD VSS sg13g2_decap_8
XFILLER_56_857 VDD VSS sg13g2_decap_8
X_1379_ _1379_/Y _1379_/A _1465_/C VDD VSS sg13g2_nand2_1
XFILLER_83_654 VDD VSS sg13g2_fill_2
XFILLER_71_805 VDD VSS sg13g2_decap_8
XFILLER_82_142 VDD VSS sg13g2_decap_8
XFILLER_83_698 VDD VSS sg13g2_decap_8
XFILLER_36_581 VDD VSS sg13g2_decap_8
XFILLER_24_721 VDD VSS sg13g2_decap_8
XFILLER_23_231 VDD VSS sg13g2_decap_8
XFILLER_51_551 VDD VSS sg13g2_decap_8
XFILLER_24_798 VDD VSS sg13g2_decap_8
XFILLER_12_938 VDD VSS sg13g2_decap_8
XFILLER_11_448 VDD VSS sg13g2_decap_8
XFILLER_23_56 VDD VSS sg13g2_decap_8
XFILLER_109_347 VDD VSS sg13g2_decap_8
XFILLER_99_49 VDD VSS sg13g2_decap_8
XIO_BOND_out_valid_pad out_valid_PAD bondpad_70x70
XFILLER_3_658 VDD VSS sg13g2_decap_8
XFILLER_79_927 VDD VSS sg13g2_fill_2
XFILLER_78_426 VDD VSS sg13g2_fill_1
XFILLER_2_168 VDD VSS sg13g2_decap_8
XFILLER_63_1060 VDD VSS sg13g2_fill_1
XFILLER_48_42 VDD VSS sg13g2_decap_8
XFILLER_24_1022 VDD VSS sg13g2_decap_8
XFILLER_59_651 VDD VSS sg13g2_decap_8
XFILLER_47_824 VDD VSS sg13g2_decap_8
XFILLER_19_504 VDD VSS sg13g2_decap_8
XFILLER_111_1036 VDD VSS sg13g2_decap_8
XFILLER_74_621 VDD VSS sg13g2_decap_4
XFILLER_74_610 VDD VSS sg13g2_fill_1
XFILLER_48_97 VDD VSS sg13g2_decap_8
XFILLER_58_161 VDD VSS sg13g2_decap_4
XFILLER_104_70 VDD VSS sg13g2_decap_8
XFILLER_58_194 VDD VSS sg13g2_decap_8
XFILLER_0_49 VDD VSS sg13g2_decap_8
XFILLER_46_367 VDD VSS sg13g2_fill_2
XFILLER_73_164 VDD VSS sg13g2_decap_8
XFILLER_27_581 VDD VSS sg13g2_decap_8
XFILLER_15_721 VDD VSS sg13g2_decap_8
XFILLER_34_518 VDD VSS sg13g2_decap_8
XFILLER_14_231 VDD VSS sg13g2_decap_8
XFILLER_70_871 VDD VSS sg13g2_decap_8
XFILLER_42_562 VDD VSS sg13g2_fill_2
XFILLER_9_14 VDD VSS sg13g2_decap_8
XFILLER_42_595 VDD VSS sg13g2_decap_8
XFILLER_30_735 VDD VSS sg13g2_decap_8
XFILLER_15_798 VDD VSS sg13g2_decap_8
XFILLER_80_84 VDD VSS sg13g2_decap_8
XFILLER_31_1015 VDD VSS sg13g2_decap_8
XFILLER_7_931 VDD VSS sg13g2_decap_8
XFILLER_6_441 VDD VSS sg13g2_decap_8
X_2351_ _2351__97/L_HI VSS VDD _2351_/D _2351_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_97_757 VDD VSS sg13g2_decap_8
X_1302_ _1302_/Y _1322_/B1 hold334/X _1322_/A2 _2345_/Q VDD VSS sg13g2_a22oi_1
XFILLER_96_245 VDD VSS sg13g2_decap_8
X_2282_ _2282_/RESET_B VSS VDD _2282_/D _2282_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_111_567 VDD VSS sg13g2_decap_8
X_1233_ _1365_/B _2355_/Q _1236_/C _1409_/C VDD VSS sg13g2_nand3_1
XFILLER_78_993 VDD VSS sg13g2_decap_8
XFILLER_38_835 VDD VSS sg13g2_decap_8
XFILLER_49_161 VDD VSS sg13g2_decap_8
XFILLER_37_301 VDD VSS sg13g2_decap_8
XFILLER_65_665 VDD VSS sg13g2_decap_4
XFILLER_80_602 VDD VSS sg13g2_decap_8
XFILLER_92_484 VDD VSS sg13g2_decap_8
XFILLER_53_838 VDD VSS sg13g2_decap_8
XFILLER_64_164 VDD VSS sg13g2_decap_8
XFILLER_25_518 VDD VSS sg13g2_decap_8
XFILLER_37_378 VDD VSS sg13g2_decap_8
XFILLER_52_359 VDD VSS sg13g2_fill_2
XFILLER_18_581 VDD VSS sg13g2_decap_8
XFILLER_100_28 VDD VSS sg13g2_decap_8
XFILLER_61_893 VDD VSS sg13g2_decap_8
XFILLER_33_595 VDD VSS sg13g2_decap_8
XFILLER_21_735 VDD VSS sg13g2_decap_8
XFILLER_60_370 VDD VSS sg13g2_fill_1
X_1997_ _1991_/X VDD _1997_/Y VSS _2071_/B _1996_/Y sg13g2_o21ai_1
XFILLER_20_245 VDD VSS sg13g2_decap_8
XFILLER_107_807 VDD VSS sg13g2_decap_8
XFILLER_87_201 VDD VSS sg13g2_decap_8
XFILLER_47_1055 VDD VSS sg13g2_decap_4
XFILLER_88_757 VDD VSS sg13g2_decap_4
XFILLER_69_971 VDD VSS sg13g2_decap_8
XFILLER_75_418 VDD VSS sg13g2_decap_8
XFILLER_28_301 VDD VSS sg13g2_decap_8
XFILLER_56_665 VDD VSS sg13g2_decap_8
XFILLER_29_868 VDD VSS sg13g2_decap_8
XFILLER_18_56 VDD VSS sg13g2_decap_8
XFILLER_83_473 VDD VSS sg13g2_decap_8
XFILLER_56_687 VDD VSS sg13g2_fill_2
XFILLER_55_175 VDD VSS sg13g2_decap_8
XFILLER_16_518 VDD VSS sg13g2_decap_8
XFILLER_28_378 VDD VSS sg13g2_decap_8
XFILLER_71_668 VDD VSS sg13g2_decap_8
XFILLER_70_112 VDD VSS sg13g2_decap_8
XFILLER_54_1004 VDD VSS sg13g2_decap_8
XFILLER_24_595 VDD VSS sg13g2_decap_8
XFILLER_51_381 VDD VSS sg13g2_decap_8
XFILLER_12_735 VDD VSS sg13g2_decap_8
XFILLER_34_77 VDD VSS sg13g2_decap_8
XFILLER_11_245 VDD VSS sg13g2_decap_8
XFILLER_8_728 VDD VSS sg13g2_decap_8
XFILLER_7_238 VDD VSS sg13g2_decap_8
XFILLER_50_21 VDD VSS sg13g2_decap_8
XFILLER_109_133 VDD VSS sg13g2_decap_8
XFILLER_50_65 VDD VSS sg13g2_decap_8
XFILLER_4_945 VDD VSS sg13g2_decap_8
XFILLER_106_895 VDD VSS sg13g2_decap_8
XFILLER_105_372 VDD VSS sg13g2_decap_8
XFILLER_3_455 VDD VSS sg13g2_decap_8
XFILLER_79_757 VDD VSS sg13g2_decap_8
XFILLER_61_1019 VDD VSS sg13g2_decap_8
XFILLER_94_727 VDD VSS sg13g2_decap_8
XFILLER_94_738 VDD VSS sg13g2_fill_1
XFILLER_93_226 VDD VSS sg13g2_decap_8
XFILLER_78_289 VDD VSS sg13g2_fill_2
XFILLER_19_301 VDD VSS sg13g2_decap_8
XFILLER_75_963 VDD VSS sg13g2_decap_8
XFILLER_35_805 VDD VSS sg13g2_decap_8
XFILLER_46_131 VDD VSS sg13g2_decap_8
XFILLER_75_996 VDD VSS sg13g2_decap_8
XFILLER_75_84 VDD VSS sg13g2_decap_8
XFILLER_62_624 VDD VSS sg13g2_decap_8
XFILLER_47_698 VDD VSS sg13g2_decap_8
XFILLER_19_378 VDD VSS sg13g2_decap_8
XFILLER_34_315 VDD VSS sg13g2_decap_8
XFILLER_90_944 VDD VSS sg13g2_fill_1
XFILLER_62_679 VDD VSS sg13g2_decap_8
XFILLER_50_819 VDD VSS sg13g2_decap_8
XFILLER_61_178 VDD VSS sg13g2_decap_8
X_1920_ _1920_/A _1920_/B _1921_/B VDD VSS sg13g2_nor2_1
XFILLER_15_595 VDD VSS sg13g2_decap_8
XFILLER_42_370 VDD VSS sg13g2_decap_8
X_1851_ _1850_/Y VDD _1852_/C VSS _1856_/A _1856_/B sg13g2_o21ai_1
XFILLER_30_532 VDD VSS sg13g2_decap_8
X_1782_ _2220_/Q _2212_/Q _1782_/Y VDD VSS sg13g2_nor2b_1
X_2342__135 VDD VSS _2342_/RESET_B sg13g2_tiehi
XFILLER_112_854 VDD VSS sg13g2_decap_8
X_2334_ _2334_/RESET_B VSS VDD _2334_/D _2334_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_58_908 VDD VSS sg13g2_decap_8
XFILLER_111_364 VDD VSS sg13g2_decap_8
XFILLER_69_267 VDD VSS sg13g2_decap_8
XFILLER_57_418 VDD VSS sg13g2_decap_8
XFILLER_27_0 VDD VSS sg13g2_decap_8
XFILLER_85_749 VDD VSS sg13g2_fill_2
XFILLER_38_632 VDD VSS sg13g2_decap_8
X_2265_ _2265_/RESET_B VSS VDD _2265_/D _2265_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_81_900 VDD VSS sg13g2_decap_8
X_1216_ VDD _1776_/A _2218_/Q VSS sg13g2_inv_1
XFILLER_84_248 VDD VSS sg13g2_decap_8
XFILLER_66_963 VDD VSS sg13g2_decap_8
X_2196_ _2196_/RESET_B VSS VDD _2196_/D _2196_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_26_805 VDD VSS sg13g2_decap_8
XFILLER_65_440 VDD VSS sg13g2_fill_1
XFILLER_92_270 VDD VSS sg13g2_decap_8
XFILLER_65_473 VDD VSS sg13g2_decap_8
XFILLER_1_70 VDD VSS sg13g2_decap_8
XFILLER_25_315 VDD VSS sg13g2_decap_8
XFILLER_37_175 VDD VSS sg13g2_decap_8
XFILLER_80_432 VDD VSS sg13g2_decap_8
XFILLER_111_49 VDD VSS sg13g2_decap_8
XFILLER_40_307 VDD VSS sg13g2_decap_8
XFILLER_52_167 VDD VSS sg13g2_decap_4
XFILLER_34_882 VDD VSS sg13g2_decap_8
XFILLER_21_532 VDD VSS sg13g2_decap_8
XFILLER_33_392 VDD VSS sg13g2_decap_8
XFILLER_101_1002 VDD VSS sg13g2_decap_4
XFILLER_107_604 VDD VSS sg13g2_decap_8
XFILLER_14_1043 VDD VSS sg13g2_decap_8
XFILLER_84_1008 VDD VSS sg13g2_decap_4
XFILLER_106_147 VDD VSS sg13g2_decap_8
XFILLER_105_7 VDD VSS sg13g2_decap_8
XFILLER_20_35 VDD VSS sg13g2_decap_8
XFILLER_88_510 VDD VSS sg13g2_decap_8
XFILLER_103_854 VDD VSS sg13g2_fill_2
XFILLER_96_28 VDD VSS sg13g2_decap_8
XFILLER_1_959 VDD VSS sg13g2_decap_8
XFILLER_88_554 VDD VSS sg13g2_decap_8
XFILLER_76_727 VDD VSS sg13g2_decap_8
XFILLER_0_469 VDD VSS sg13g2_decap_8
XFILLER_69_790 VDD VSS sg13g2_decap_8
XFILLER_102_375 VDD VSS sg13g2_decap_8
XFILLER_75_215 VDD VSS sg13g2_decap_8
XFILLER_29_77 VDD VSS sg13g2_decap_8
XFILLER_21_1036 VDD VSS sg13g2_decap_8
XFILLER_29_665 VDD VSS sg13g2_decap_8
XFILLER_56_440 VDD VSS sg13g2_decap_8
XFILLER_17_805 VDD VSS sg13g2_decap_8
XFILLER_44_613 VDD VSS sg13g2_decap_8
XFILLER_16_315 VDD VSS sg13g2_decap_8
XFILLER_45_21 VDD VSS sg13g2_decap_8
XFILLER_28_175 VDD VSS sg13g2_decap_8
XFILLER_72_955 VDD VSS sg13g2_decap_8
XFILLER_83_292 VDD VSS sg13g2_decap_8
XFILLER_71_432 VDD VSS sg13g2_decap_8
XFILLER_43_112 VDD VSS sg13g2_decap_8
XFILLER_32_819 VDD VSS sg13g2_decap_8
XFILLER_43_156 VDD VSS sg13g2_fill_1
XFILLER_40_830 VDD VSS sg13g2_decap_8
XFILLER_25_882 VDD VSS sg13g2_decap_8
XFILLER_31_329 VDD VSS sg13g2_decap_8
XFILLER_43_189 VDD VSS sg13g2_decap_8
XFILLER_12_532 VDD VSS sg13g2_decap_8
XFILLER_61_42 VDD VSS sg13g2_decap_8
XFILLER_24_392 VDD VSS sg13g2_decap_8
XFILLER_8_525 VDD VSS sg13g2_decap_8
XFILLER_61_97 VDD VSS sg13g2_fill_2
XFILLER_99_808 VDD VSS sg13g2_fill_2
Xin_ready_pad _2355_/Q IOVDD IOVSS in_ready_PAD VDD VSS sg13g2_IOPadOut30mA
XFILLER_4_742 VDD VSS sg13g2_decap_8
XFILLER_98_318 VDD VSS sg13g2_decap_8
XFILLER_3_252 VDD VSS sg13g2_decap_8
XFILLER_106_692 VDD VSS sg13g2_decap_8
XFILLER_79_554 VDD VSS sg13g2_decap_8
XFILLER_67_705 VDD VSS sg13g2_fill_2
XFILLER_6_1008 VDD VSS sg13g2_decap_8
XFILLER_48_930 VDD VSS sg13g2_decap_8
XFILLER_20_7 VDD VSS sg13g2_decap_8
XFILLER_39_429 VDD VSS sg13g2_decap_8
X_2050_ _1922_/Y _1953_/A _2069_/S _2050_/X VDD VSS sg13g2_mux2_1
XFILLER_75_782 VDD VSS sg13g2_decap_8
XFILLER_48_974 VDD VSS sg13g2_decap_8
XFILLER_35_602 VDD VSS sg13g2_decap_8
XFILLER_47_451 VDD VSS sg13g2_decap_4
XFILLER_62_421 VDD VSS sg13g2_decap_8
XFILLER_19_175 VDD VSS sg13g2_decap_8
XFILLER_34_112 VDD VSS sg13g2_decap_8
XFILLER_47_495 VDD VSS sg13g2_decap_8
XFILLER_90_752 VDD VSS sg13g2_decap_8
XFILLER_35_679 VDD VSS sg13g2_decap_8
XFILLER_23_819 VDD VSS sg13g2_decap_8
XFILLER_37_1043 VDD VSS sg13g2_decap_8
XFILLER_62_498 VDD VSS sg13g2_fill_2
XFILLER_16_882 VDD VSS sg13g2_decap_8
XFILLER_22_329 VDD VSS sg13g2_decap_8
XFILLER_34_189 VDD VSS sg13g2_decap_8
X_1903_ _1903_/B _1903_/A _1943_/A VDD VSS sg13g2_xor2_1
XFILLER_15_392 VDD VSS sg13g2_decap_8
XFILLER_31_896 VDD VSS sg13g2_decap_8
X_1834_ _2246_/Q _2205_/Q _1920_/A VDD VSS sg13g2_nor2b_1
XIO_FILL_IO_SOUTH_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_1765_ _1766_/B _1926_/B _1940_/A VDD VSS sg13g2_nand2_1
Xhold514 _2317_/Q VDD VSS hold514/X sg13g2_dlygate4sd3_1
Xhold525 _2226_/Q VDD VSS hold525/X sg13g2_dlygate4sd3_1
Xhold536 _2242_/Q VDD VSS hold536/X sg13g2_dlygate4sd3_1
Xhold503 _2314_/Q VDD VSS hold503/X sg13g2_dlygate4sd3_1
XFILLER_89_307 VDD VSS sg13g2_decap_8
X_1696_ _1725_/A _1696_/B _1696_/Y VDD VSS sg13g2_nor2_1
Xhold558 _1258_/Y VDD VSS _2356_/D sg13g2_dlygate4sd3_1
Xhold569 _2355_/Q VDD VSS hold569/X sg13g2_dlygate4sd3_1
Xhold547 _2292_/Q VDD VSS hold547/X sg13g2_dlygate4sd3_1
XFILLER_83_1052 VDD VSS sg13g2_decap_8
XFILLER_98_841 VDD VSS sg13g2_decap_8
XFILLER_112_651 VDD VSS sg13g2_decap_8
XFILLER_106_49 VDD VSS sg13g2_decap_8
X_2317_ _2317_/RESET_B VSS VDD _2317_/D _2317_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_111_161 VDD VSS sg13g2_decap_8
X_2320__230 VDD VSS _2320_/RESET_B sg13g2_tiehi
XFILLER_44_1047 VDD VSS sg13g2_decap_8
XFILLER_58_749 VDD VSS sg13g2_decap_4
XFILLER_100_868 VDD VSS sg13g2_decap_8
XFILLER_85_568 VDD VSS sg13g2_decap_8
XFILLER_39_941 VDD VSS sg13g2_decap_8
X_2248_ _2248_/RESET_B VSS VDD _2248_/D _2248_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_72_207 VDD VSS sg13g2_decap_8
XFILLER_66_782 VDD VSS sg13g2_fill_2
XFILLER_26_602 VDD VSS sg13g2_decap_8
XFILLER_54_955 VDD VSS sg13g2_decap_8
X_2179_ _2179_/RESET_B VSS VDD _2179_/D _2179_/Q _2365_/CLK sg13g2_dfrbpq_1
X_2277__195 VDD VSS _2277_/RESET_B sg13g2_tiehi
XFILLER_53_410 VDD VSS sg13g2_decap_4
XFILLER_25_112 VDD VSS sg13g2_decap_8
XFILLER_38_495 VDD VSS sg13g2_decap_8
XFILLER_26_679 VDD VSS sg13g2_decap_8
XFILLER_14_819 VDD VSS sg13g2_decap_8
XFILLER_90_1001 VDD VSS sg13g2_decap_8
XFILLER_80_262 VDD VSS sg13g2_decap_8
XFILLER_53_498 VDD VSS sg13g2_decap_8
XFILLER_13_329 VDD VSS sg13g2_decap_8
XFILLER_15_35 VDD VSS sg13g2_decap_8
XFILLER_40_126 VDD VSS sg13g2_decap_8
XFILLER_25_189 VDD VSS sg13g2_decap_8
XFILLER_22_896 VDD VSS sg13g2_decap_8
XFILLER_108_913 VDD VSS sg13g2_decap_8
XFILLER_31_56 VDD VSS sg13g2_decap_8
XFILLER_107_423 VDD VSS sg13g2_decap_8
XFILLER_5_539 VDD VSS sg13g2_decap_8
XFILLER_103_651 VDD VSS sg13g2_decap_8
XFILLER_89_852 VDD VSS sg13g2_decap_8
XFILLER_1_756 VDD VSS sg13g2_decap_8
XFILLER_88_373 VDD VSS sg13g2_decap_8
XFILLER_102_161 VDD VSS sg13g2_decap_8
XFILLER_0_266 VDD VSS sg13g2_decap_8
XFILLER_76_557 VDD VSS sg13g2_decap_8
XFILLER_48_237 VDD VSS sg13g2_decap_8
XFILLER_48_248 VDD VSS sg13g2_fill_1
XFILLER_17_602 VDD VSS sg13g2_decap_8
XFILLER_29_462 VDD VSS sg13g2_decap_8
XFILLER_91_549 VDD VSS sg13g2_decap_8
XFILLER_45_933 VDD VSS sg13g2_decap_8
XFILLER_57_793 VDD VSS sg13g2_decap_8
XFILLER_56_270 VDD VSS sg13g2_decap_8
XFILLER_16_112 VDD VSS sg13g2_decap_8
XFILLER_44_432 VDD VSS sg13g2_decap_8
XFILLER_112_70 VDD VSS sg13g2_decap_8
XFILLER_60_914 VDD VSS sg13g2_decap_8
XFILLER_17_679 VDD VSS sg13g2_decap_8
XFILLER_32_616 VDD VSS sg13g2_decap_8
XFILLER_16_189 VDD VSS sg13g2_decap_8
XFILLER_44_476 VDD VSS sg13g2_fill_1
XFILLER_72_63 VDD VSS sg13g2_decap_8
XFILLER_31_126 VDD VSS sg13g2_decap_8
XFILLER_9_812 VDD VSS sg13g2_decap_8
XFILLER_13_896 VDD VSS sg13g2_decap_8
XFILLER_8_322 VDD VSS sg13g2_decap_8
XFILLER_9_889 VDD VSS sg13g2_decap_8
XFILLER_68_7 VDD VSS sg13g2_decap_8
X_1550_ VDD _1550_/Y _1550_/A VSS sg13g2_inv_1
XFILLER_8_399 VDD VSS sg13g2_decap_8
XFILLER_67_1025 VDD VSS sg13g2_decap_8
XFILLER_98_126 VDD VSS sg13g2_decap_8
X_1481_ VSS VDD _1194_/Y _1481_/A2 _2259_/D _1480_/Y sg13g2_a21oi_1
XFILLER_95_822 VDD VSS sg13g2_decap_8
XFILLER_94_310 VDD VSS sg13g2_decap_8
XFILLER_79_384 VDD VSS sg13g2_decap_8
XFILLER_67_546 VDD VSS sg13g2_decap_8
XFILLER_39_259 VDD VSS sg13g2_decap_8
X_2102_ _2102_/B _2102_/C _2102_/A _2104_/B VDD VSS sg13g2_nand3_1
XFILLER_94_354 VDD VSS sg13g2_fill_2
XFILLER_82_527 VDD VSS sg13g2_decap_8
XFILLER_48_782 VDD VSS sg13g2_decap_8
X_2033_ _2034_/B _2033_/B _2004_/B VDD VSS sg13g2_nand2b_1
XFILLER_94_398 VDD VSS sg13g2_decap_8
XFILLER_63_730 VDD VSS sg13g2_decap_8
XFILLER_48_793 VDD VSS sg13g2_decap_8
XFILLER_47_292 VDD VSS sg13g2_decap_8
XFILLER_36_966 VDD VSS sg13g2_decap_8
XFILLER_51_925 VDD VSS sg13g2_decap_8
XFILLER_23_616 VDD VSS sg13g2_decap_8
XFILLER_62_273 VDD VSS sg13g2_decap_8
XFILLER_35_476 VDD VSS sg13g2_decap_8
XFILLER_50_402 VDD VSS sg13g2_decap_8
XFILLER_94_0 VDD VSS sg13g2_decap_8
XFILLER_22_126 VDD VSS sg13g2_decap_8
XFILLER_50_479 VDD VSS sg13g2_decap_8
XFILLER_31_693 VDD VSS sg13g2_decap_8
X_1817_ _1819_/B _1929_/B _1817_/B _1939_/B VDD VSS sg13g2_and3_1
Xhold311 _1286_/Y VDD VSS _1287_/A sg13g2_dlygate4sd3_1
XFILLER_7_91 VDD VSS sg13g2_decap_8
Xhold300 _2108_/Y VDD VSS _2354_/D sg13g2_dlygate4sd3_1
Xhold322 _2167_/Q VDD VSS hold322/X sg13g2_dlygate4sd3_1
Xhold344 _1324_/Y VDD VSS _1325_/A sg13g2_dlygate4sd3_1
Xhold333 _1296_/Y VDD VSS _1297_/A sg13g2_dlygate4sd3_1
X_1748_ _1751_/B _2240_/Q _2232_/Q VDD VSS sg13g2_nand2b_1
XFILLER_11_1057 VDD VSS sg13g2_decap_4
XFILLER_105_938 VDD VSS sg13g2_decap_8
Xhold355 _2174_/Q VDD VSS hold355/X sg13g2_dlygate4sd3_1
Xhold366 _2200_/Q VDD VSS hold366/X sg13g2_dlygate4sd3_1
Xhold377 _2189_/Q VDD VSS hold377/X sg13g2_dlygate4sd3_1
XFILLER_104_437 VDD VSS sg13g2_decap_8
XFILLER_89_126 VDD VSS sg13g2_decap_8
X_1679_ _1680_/B _1679_/B _2311_/D VDD VSS sg13g2_and2_1
Xhold388 _1306_/Y VDD VSS _1307_/A sg13g2_dlygate4sd3_1
Xhold399 _2199_/Q VDD VSS hold399/X sg13g2_dlygate4sd3_1
XFILLER_86_855 VDD VSS sg13g2_decap_8
XFILLER_85_376 VDD VSS sg13g2_decap_8
XFILLER_73_505 VDD VSS sg13g2_decap_4
XFILLER_58_579 VDD VSS sg13g2_fill_1
XFILLER_46_719 VDD VSS sg13g2_decap_8
XFILLER_73_538 VDD VSS sg13g2_decap_8
XFILLER_27_966 VDD VSS sg13g2_decap_8
XFILLER_42_903 VDD VSS sg13g2_decap_8
XFILLER_26_56 VDD VSS sg13g2_decap_8
XFILLER_14_616 VDD VSS sg13g2_decap_8
XFILLER_26_476 VDD VSS sg13g2_decap_8
XFILLER_41_402 VDD VSS sg13g2_decap_8
XFILLER_13_126 VDD VSS sg13g2_decap_8
XFILLER_107_1052 VDD VSS sg13g2_decap_8
X_2212__116 VDD VSS _2212_/RESET_B sg13g2_tiehi
XFILLER_9_119 VDD VSS sg13g2_decap_8
XFILLER_22_693 VDD VSS sg13g2_decap_8
XFILLER_10_833 VDD VSS sg13g2_decap_8
XFILLER_42_77 VDD VSS sg13g2_decap_8
XFILLER_108_710 VDD VSS sg13g2_decap_8
XFILLER_6_826 VDD VSS sg13g2_decap_8
XFILLER_5_336 VDD VSS sg13g2_decap_8
XFILLER_108_787 VDD VSS sg13g2_decap_8
XFILLER_1_553 VDD VSS sg13g2_decap_8
XFILLER_104_971 VDD VSS sg13g2_decap_8
XFILLER_89_671 VDD VSS sg13g2_decap_8
XFILLER_107_70 VDD VSS sg13g2_decap_8
X_2309__79 VDD VSS _2309__79/L_HI sg13g2_tiehi
XFILLER_3_49 VDD VSS sg13g2_decap_8
XFILLER_77_844 VDD VSS sg13g2_decap_8
XFILLER_67_63 VDD VSS sg13g2_decap_8
XFILLER_77_877 VDD VSS sg13g2_decap_8
XFILLER_49_579 VDD VSS sg13g2_decap_8
XFILLER_92_847 VDD VSS sg13g2_decap_8
XFILLER_76_387 VDD VSS sg13g2_decap_8
XFILLER_57_590 VDD VSS sg13g2_fill_1
XFILLER_91_368 VDD VSS sg13g2_decap_8
XFILLER_33_903 VDD VSS sg13g2_decap_8
XFILLER_18_966 VDD VSS sg13g2_decap_8
XFILLER_83_84 VDD VSS sg13g2_decap_8
XFILLER_60_722 VDD VSS sg13g2_decap_8
XFILLER_17_476 VDD VSS sg13g2_decap_8
XFILLER_32_413 VDD VSS sg13g2_decap_8
XFILLER_60_755 VDD VSS sg13g2_decap_8
XFILLER_73_1051 VDD VSS sg13g2_decap_8
XFILLER_60_799 VDD VSS sg13g2_decap_8
XFILLER_34_1057 VDD VSS sg13g2_decap_4
XFILLER_13_693 VDD VSS sg13g2_decap_8
XFILLER_9_686 VDD VSS sg13g2_decap_8
XFILLER_8_196 VDD VSS sg13g2_decap_8
X_1602_ _1639_/A _1602_/B hold562/X VDD VSS sg13g2_nand2b_1
XFILLER_99_435 VDD VSS sg13g2_decap_8
X_1533_ _1534_/B _1527_/Y _1532_/Y hold520/X _1527_/B VDD VSS sg13g2_a22oi_1
X_1464_ VSS VDD _1388_/Y _1455_/B _2251_/D _1463_/Y sg13g2_a21oi_1
XFILLER_80_1033 VDD VSS sg13g2_fill_1
XFILLER_101_407 VDD VSS sg13g2_decap_4
XFILLER_95_630 VDD VSS sg13g2_decap_8
X_1395_ _1396_/A _1392_/Y hold554/X _1392_/B _1370_/A VDD VSS sg13g2_a22oi_1
XFILLER_41_1028 VDD VSS sg13g2_decap_8
XFILLER_68_855 VDD VSS sg13g2_decap_8
XFILLER_67_343 VDD VSS sg13g2_decap_8
XFILLER_110_963 VDD VSS sg13g2_decap_8
XFILLER_94_140 VDD VSS sg13g2_decap_8
XFILLER_67_376 VDD VSS sg13g2_fill_1
XFILLER_83_836 VDD VSS sg13g2_fill_2
XFILLER_82_335 VDD VSS sg13g2_decap_8
XFILLER_82_313 VDD VSS sg13g2_fill_2
XFILLER_103_28 VDD VSS sg13g2_decap_8
X_2016_ _2021_/S _1901_/B _1914_/A _1949_/A _1889_/A _2022_/S _2017_/B VDD VSS sg13g2_mux4_1
XFILLER_82_368 VDD VSS sg13g2_fill_2
XFILLER_36_763 VDD VSS sg13g2_decap_8
XFILLER_24_903 VDD VSS sg13g2_decap_8
XFILLER_23_413 VDD VSS sg13g2_decap_8
XFILLER_35_273 VDD VSS sg13g2_decap_8
XFILLER_51_744 VDD VSS sg13g2_decap_8
XFILLER_32_980 VDD VSS sg13g2_decap_8
XFILLER_109_518 VDD VSS sg13g2_decap_8
XFILLER_12_14 VDD VSS sg13g2_decap_8
XFILLER_31_490 VDD VSS sg13g2_decap_8
XFILLER_105_735 VDD VSS sg13g2_decap_8
XFILLER_104_245 VDD VSS sg13g2_decap_8
XFILLER_86_630 VDD VSS sg13g2_decap_8
XFILLER_98_490 VDD VSS sg13g2_decap_8
XFILLER_59_844 VDD VSS sg13g2_decap_4
XFILLER_101_963 VDD VSS sg13g2_decap_8
XFILLER_74_814 VDD VSS sg13g2_decap_8
XFILLER_58_365 VDD VSS sg13g2_decap_8
XFILLER_58_376 VDD VSS sg13g2_fill_1
XFILLER_100_484 VDD VSS sg13g2_decap_8
XFILLER_2_1022 VDD VSS sg13g2_decap_8
XFILLER_74_869 VDD VSS sg13g2_decap_4
XIO_BOND_out_data_pads\[3\].out_data_pad out_data_PADs[3] bondpad_70x70
XFILLER_27_763 VDD VSS sg13g2_decap_8
XFILLER_15_903 VDD VSS sg13g2_decap_8
XFILLER_37_77 VDD VSS sg13g2_decap_8
XFILLER_73_379 VDD VSS sg13g2_decap_8
XFILLER_57_1024 VDD VSS sg13g2_decap_8
XFILLER_57_1035 VDD VSS sg13g2_fill_2
XFILLER_54_582 VDD VSS sg13g2_decap_8
XFILLER_42_700 VDD VSS sg13g2_decap_8
XFILLER_14_413 VDD VSS sg13g2_decap_8
XFILLER_26_273 VDD VSS sg13g2_decap_8
XFILLER_57_1046 VDD VSS sg13g2_decap_8
XFILLER_54_593 VDD VSS sg13g2_fill_1
XFILLER_18_1008 VDD VSS sg13g2_decap_8
XFILLER_30_917 VDD VSS sg13g2_decap_8
XFILLER_42_777 VDD VSS sg13g2_decap_8
XFILLER_53_87 VDD VSS sg13g2_fill_2
XFILLER_53_76 VDD VSS sg13g2_decap_8
XFILLER_23_980 VDD VSS sg13g2_decap_8
XFILLER_41_287 VDD VSS sg13g2_decap_8
XFILLER_10_630 VDD VSS sg13g2_decap_8
XFILLER_22_490 VDD VSS sg13g2_decap_8
XFILLER_6_623 VDD VSS sg13g2_decap_8
XFILLER_5_133 VDD VSS sg13g2_decap_8
XFILLER_108_584 VDD VSS sg13g2_decap_8
XFILLER_64_1028 VDD VSS sg13g2_decap_8
XFILLER_2_840 VDD VSS sg13g2_decap_8
XFILLER_96_427 VDD VSS sg13g2_decap_8
XFILLER_78_84 VDD VSS sg13g2_decap_8
XFILLER_1_350 VDD VSS sg13g2_decap_8
XFILLER_111_749 VDD VSS sg13g2_decap_8
XFILLER_77_674 VDD VSS sg13g2_decap_8
XFILLER_110_259 VDD VSS sg13g2_decap_8
XFILLER_76_140 VDD VSS sg13g2_decap_8
X_2297__121 VDD VSS _2297_/RESET_B sg13g2_tiehi
XFILLER_64_335 VDD VSS sg13g2_decap_4
XFILLER_49_398 VDD VSS sg13g2_decap_8
X_2338__151 VDD VSS _2338_/RESET_B sg13g2_tiehi
XFILLER_18_763 VDD VSS sg13g2_decap_8
XFILLER_80_839 VDD VSS sg13g2_decap_8
XFILLER_45_560 VDD VSS sg13g2_decap_8
XFILLER_33_700 VDD VSS sg13g2_decap_8
XFILLER_52_519 VDD VSS sg13g2_decap_8
XFILLER_17_273 VDD VSS sg13g2_decap_8
XFILLER_32_210 VDD VSS sg13g2_decap_8
XFILLER_21_917 VDD VSS sg13g2_decap_8
XFILLER_60_552 VDD VSS sg13g2_decap_8
XFILLER_33_777 VDD VSS sg13g2_decap_8
XFILLER_20_427 VDD VSS sg13g2_decap_8
XFILLER_14_980 VDD VSS sg13g2_decap_8
XFILLER_32_287 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_12_clk clkbuf_2_2__f_clk/X clkload9/A VDD VSS sg13g2_buf_8
XFILLER_13_490 VDD VSS sg13g2_decap_8
XFILLER_9_483 VDD VSS sg13g2_decap_8
X_2165__210 VDD VSS _2165_/RESET_B sg13g2_tiehi
XFILLER_57_0 VDD VSS sg13g2_decap_8
XFILLER_99_221 VDD VSS sg13g2_decap_8
X_1516_ VSS VDD _1516_/X _1516_/B _1516_/A sg13g2_or2_1
XFILLER_88_928 VDD VSS sg13g2_fill_1
XFILLER_87_416 VDD VSS sg13g2_decap_8
XFILLER_4_70 VDD VSS sg13g2_decap_8
XFILLER_101_248 VDD VSS sg13g2_decap_8
X_1447_ _1492_/A _1495_/C _1493_/A VDD VSS sg13g2_and2_1
XFILLER_96_961 VDD VSS sg13g2_fill_2
XFILLER_110_760 VDD VSS sg13g2_decap_8
X_1378_ _1377_/Y VDD _2214_/D VSS _1367_/B _1376_/Y sg13g2_o21ai_1
XFILLER_68_652 VDD VSS sg13g2_decap_8
XFILLER_83_633 VDD VSS sg13g2_decap_8
XFILLER_83_677 VDD VSS sg13g2_decap_8
XFILLER_67_195 VDD VSS sg13g2_decap_8
XFILLER_55_368 VDD VSS sg13g2_decap_4
XFILLER_70_327 VDD VSS sg13g2_decap_4
XFILLER_64_880 VDD VSS sg13g2_decap_8
XFILLER_36_560 VDD VSS sg13g2_decap_8
XFILLER_24_700 VDD VSS sg13g2_decap_8
XFILLER_55_379 VDD VSS sg13g2_fill_1
XFILLER_51_530 VDD VSS sg13g2_decap_8
XFILLER_23_210 VDD VSS sg13g2_decap_8
XFILLER_24_777 VDD VSS sg13g2_decap_8
XFILLER_12_917 VDD VSS sg13g2_decap_8
XFILLER_11_427 VDD VSS sg13g2_decap_8
XFILLER_23_35 VDD VSS sg13g2_decap_8
XFILLER_23_287 VDD VSS sg13g2_decap_8
XFILLER_104_1055 VDD VSS sg13g2_decap_4
XFILLER_99_28 VDD VSS sg13g2_decap_8
XFILLER_20_994 VDD VSS sg13g2_decap_8
XFILLER_3_637 VDD VSS sg13g2_decap_8
XFILLER_2_147 VDD VSS sg13g2_decap_8
XFILLER_24_1001 VDD VSS sg13g2_decap_8
XFILLER_59_630 VDD VSS sg13g2_decap_8
XFILLER_48_21 VDD VSS sg13g2_decap_8
XFILLER_87_972 VDD VSS sg13g2_fill_2
XFILLER_87_983 VDD VSS sg13g2_decap_8
XFILLER_111_1015 VDD VSS sg13g2_decap_8
XFILLER_101_793 VDD VSS sg13g2_decap_8
XFILLER_86_482 VDD VSS sg13g2_decap_8
XFILLER_59_685 VDD VSS sg13g2_decap_8
XFILLER_73_143 VDD VSS sg13g2_decap_8
XFILLER_0_28 VDD VSS sg13g2_decap_8
XFILLER_74_688 VDD VSS sg13g2_decap_8
XFILLER_27_560 VDD VSS sg13g2_decap_8
XFILLER_61_305 VDD VSS sg13g2_decap_8
XFILLER_15_700 VDD VSS sg13g2_decap_8
XFILLER_64_42 VDD VSS sg13g2_decap_8
XFILLER_46_379 VDD VSS sg13g2_decap_8
XFILLER_54_390 VDD VSS sg13g2_fill_2
XFILLER_14_210 VDD VSS sg13g2_decap_8
XFILLER_70_850 VDD VSS sg13g2_decap_8
XFILLER_42_574 VDD VSS sg13g2_decap_8
XFILLER_30_714 VDD VSS sg13g2_decap_8
XFILLER_15_777 VDD VSS sg13g2_decap_8
XFILLER_14_287 VDD VSS sg13g2_decap_8
XFILLER_80_63 VDD VSS sg13g2_decap_8
XFILLER_7_910 VDD VSS sg13g2_decap_8
Xin_data_pads\[1\].in_data_pad IOVDD IOVSS _1370_/A in_data_PADs[1] VDD VSS sg13g2_IOPadIn
XFILLER_6_420 VDD VSS sg13g2_decap_8
XFILLER_11_994 VDD VSS sg13g2_decap_8
XFILLER_109_882 VDD VSS sg13g2_decap_8
XFILLER_108_370 VDD VSS sg13g2_fill_2
XFILLER_7_987 VDD VSS sg13g2_decap_8
XFILLER_50_7 VDD VSS sg13g2_decap_8
XFILLER_6_497 VDD VSS sg13g2_decap_8
XFILLER_69_416 VDD VSS sg13g2_fill_1
X_2350_ _2350_/RESET_B VSS VDD _2350_/D _2350_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_111_546 VDD VSS sg13g2_decap_8
XFILLER_96_224 VDD VSS sg13g2_decap_8
XFILLER_69_438 VDD VSS sg13g2_fill_1
X_1301_ VDD _2180_/D _1301_/A VSS sg13g2_inv_1
X_2281_ _2281_/RESET_B VSS VDD _2281_/D _2281_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_78_972 VDD VSS sg13g2_decap_8
XFILLER_38_814 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_1_clk clkbuf_leaf_5_clk/A clkload4/A VDD VSS sg13g2_buf_8
X_1232_ _1583_/A _1234_/B _1388_/B VDD VSS sg13g2_nor2_1
XFILLER_49_140 VDD VSS sg13g2_decap_8
XFILLER_77_493 VDD VSS sg13g2_fill_1
XFILLER_77_482 VDD VSS sg13g2_decap_8
XFILLER_92_441 VDD VSS sg13g2_decap_8
XFILLER_64_143 VDD VSS sg13g2_decap_8
XFILLER_37_357 VDD VSS sg13g2_decap_8
XFILLER_93_997 VDD VSS sg13g2_decap_8
XFILLER_53_817 VDD VSS sg13g2_decap_8
XFILLER_46_880 VDD VSS sg13g2_decap_8
XFILLER_18_560 VDD VSS sg13g2_decap_8
XFILLER_61_872 VDD VSS sg13g2_decap_8
XFILLER_21_714 VDD VSS sg13g2_decap_8
XFILLER_33_574 VDD VSS sg13g2_decap_8
XFILLER_20_224 VDD VSS sg13g2_decap_8
X_1996_ _1996_/Y _1976_/Y _1995_/X _1974_/X _1973_/Y VDD VSS sg13g2_a22oi_1
XFILLER_9_280 VDD VSS sg13g2_decap_8
XFILLER_109_49 VDD VSS sg13g2_decap_8
XFILLER_88_714 VDD VSS sg13g2_decap_8
XFILLER_47_1034 VDD VSS sg13g2_decap_8
XFILLER_88_736 VDD VSS sg13g2_decap_8
XFILLER_102_535 VDD VSS sg13g2_decap_8
XFILLER_69_950 VDD VSS sg13g2_decap_8
XFILLER_29_847 VDD VSS sg13g2_decap_8
XFILLER_18_35 VDD VSS sg13g2_decap_8
XFILLER_83_452 VDD VSS sg13g2_fill_2
XFILLER_56_644 VDD VSS sg13g2_decap_8
XFILLER_28_357 VDD VSS sg13g2_decap_8
XFILLER_55_154 VDD VSS sg13g2_decap_8
XFILLER_71_647 VDD VSS sg13g2_decap_8
XFILLER_70_168 VDD VSS sg13g2_decap_8
XFILLER_24_574 VDD VSS sg13g2_decap_8
XFILLER_12_714 VDD VSS sg13g2_decap_8
XFILLER_34_56 VDD VSS sg13g2_decap_8
XFILLER_11_224 VDD VSS sg13g2_decap_8
XFILLER_8_707 VDD VSS sg13g2_decap_8
XFILLER_109_112 VDD VSS sg13g2_decap_8
XFILLER_7_217 VDD VSS sg13g2_decap_8
Xclkload0 clkload0/Y clkload0/A VDD VSS sg13g2_inv_2
XFILLER_20_791 VDD VSS sg13g2_decap_8
XFILLER_50_44 VDD VSS sg13g2_decap_8
XFILLER_109_189 VDD VSS sg13g2_decap_8
XFILLER_4_924 VDD VSS sg13g2_decap_8
XFILLER_50_99 VDD VSS sg13g2_decap_8
XFILLER_3_434 VDD VSS sg13g2_decap_8
XFILLER_106_874 VDD VSS sg13g2_decap_8
XFILLER_79_703 VDD VSS sg13g2_fill_1
XFILLER_105_351 VDD VSS sg13g2_decap_8
XFILLER_79_736 VDD VSS sg13g2_decap_8
XFILLER_59_86 VDD VSS sg13g2_fill_1
XFILLER_59_75 VDD VSS sg13g2_decap_8
XFILLER_94_706 VDD VSS sg13g2_decap_8
XFILLER_78_246 VDD VSS sg13g2_decap_8
XFILLER_8_1050 VDD VSS sg13g2_decap_8
XFILLER_87_780 VDD VSS sg13g2_decap_8
XFILLER_93_205 VDD VSS sg13g2_fill_2
XFILLER_75_63 VDD VSS sg13g2_decap_8
XFILLER_47_644 VDD VSS sg13g2_decap_8
XFILLER_19_357 VDD VSS sg13g2_decap_8
X_2259__233 VDD VSS _2259_/RESET_B sg13g2_tiehi
XFILLER_90_923 VDD VSS sg13g2_decap_8
XFILLER_62_603 VDD VSS sg13g2_decap_8
XFILLER_47_677 VDD VSS sg13g2_decap_8
XFILLER_62_669 VDD VSS sg13g2_fill_1
XFILLER_61_157 VDD VSS sg13g2_decap_8
XFILLER_98_7 VDD VSS sg13g2_decap_8
XFILLER_91_84 VDD VSS sg13g2_decap_8
XFILLER_15_574 VDD VSS sg13g2_decap_8
XFILLER_30_511 VDD VSS sg13g2_decap_8
X_1850_ _1862_/A _1850_/B _1850_/Y VDD VSS sg13g2_nor2_1
X_1781_ _2219_/Q _2211_/Q _1929_/A VDD VSS sg13g2_nor2b_1
XFILLER_30_588 VDD VSS sg13g2_decap_8
XFILLER_11_791 VDD VSS sg13g2_decap_8
XFILLER_7_784 VDD VSS sg13g2_decap_8
XFILLER_6_294 VDD VSS sg13g2_decap_8
XFILLER_112_833 VDD VSS sg13g2_decap_8
X_2333_ _2333_/RESET_B VSS VDD _2333_/D _2333_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_97_577 VDD VSS sg13g2_decap_8
XFILLER_111_343 VDD VSS sg13g2_decap_8
XFILLER_69_246 VDD VSS sg13g2_decap_8
XFILLER_85_728 VDD VSS sg13g2_decap_8
XFILLER_84_227 VDD VSS sg13g2_decap_8
XFILLER_38_611 VDD VSS sg13g2_decap_8
X_2264_ _2264_/RESET_B VSS VDD _2264_/D _2264_/Q _2365_/CLK sg13g2_dfrbpq_1
X_1215_ VDD _1215_/Y _2244_/Q VSS sg13g2_inv_1
XFILLER_66_942 VDD VSS sg13g2_decap_8
X_2195_ _2195_/RESET_B VSS VDD _2195_/D _2195_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_38_688 VDD VSS sg13g2_decap_8
XFILLER_65_452 VDD VSS sg13g2_decap_8
XFILLER_37_154 VDD VSS sg13g2_decap_8
XFILLER_81_967 VDD VSS sg13g2_decap_8
XFILLER_77_1049 VDD VSS sg13g2_decap_8
XFILLER_93_794 VDD VSS sg13g2_decap_4
XFILLER_80_411 VDD VSS sg13g2_decap_8
XFILLER_111_28 VDD VSS sg13g2_decap_8
XFILLER_52_124 VDD VSS sg13g2_decap_8
XFILLER_34_861 VDD VSS sg13g2_decap_8
XFILLER_80_488 VDD VSS sg13g2_decap_8
XFILLER_21_511 VDD VSS sg13g2_decap_8
XFILLER_33_371 VDD VSS sg13g2_decap_8
XFILLER_21_588 VDD VSS sg13g2_decap_8
XFILLER_14_1022 VDD VSS sg13g2_decap_8
X_1979_ _1978_/C VDD _1980_/B VSS _1978_/A _1978_/B sg13g2_o21ai_1
XFILLER_20_14 VDD VSS sg13g2_decap_8
XFILLER_106_126 VDD VSS sg13g2_decap_8
XFILLER_1_938 VDD VSS sg13g2_decap_8
XFILLER_103_866 VDD VSS sg13g2_fill_1
XFILLER_76_706 VDD VSS sg13g2_decap_8
XFILLER_102_354 VDD VSS sg13g2_decap_8
XFILLER_0_448 VDD VSS sg13g2_decap_8
XFILLER_29_56 VDD VSS sg13g2_decap_8
XFILLER_60_1053 VDD VSS sg13g2_decap_8
XFILLER_21_1015 VDD VSS sg13g2_decap_8
XFILLER_29_644 VDD VSS sg13g2_decap_8
XFILLER_72_912 VDD VSS sg13g2_decap_4
XFILLER_57_986 VDD VSS sg13g2_decap_8
XFILLER_28_154 VDD VSS sg13g2_decap_8
XFILLER_71_411 VDD VSS sg13g2_decap_8
XFILLER_25_861 VDD VSS sg13g2_decap_8
XFILLER_45_77 VDD VSS sg13g2_decap_8
XFILLER_31_308 VDD VSS sg13g2_decap_8
XFILLER_71_488 VDD VSS sg13g2_decap_8
XFILLER_12_511 VDD VSS sg13g2_decap_8
XFILLER_24_371 VDD VSS sg13g2_decap_8
XFILLER_52_691 VDD VSS sg13g2_decap_8
XFILLER_8_504 VDD VSS sg13g2_decap_8
XFILLER_61_21 VDD VSS sg13g2_decap_8
XFILLER_40_886 VDD VSS sg13g2_decap_8
XFILLER_12_588 VDD VSS sg13g2_decap_8
XFILLER_6_49 VDD VSS sg13g2_decap_8
XFILLER_4_721 VDD VSS sg13g2_decap_8
XFILLER_3_231 VDD VSS sg13g2_decap_8
XFILLER_106_671 VDD VSS sg13g2_decap_8
XFILLER_79_533 VDD VSS sg13g2_decap_8
XFILLER_10_91 VDD VSS sg13g2_decap_8
XFILLER_4_798 VDD VSS sg13g2_decap_8
XFILLER_79_577 VDD VSS sg13g2_decap_8
XFILLER_39_408 VDD VSS sg13g2_decap_8
XFILLER_94_503 VDD VSS sg13g2_decap_4
XFILLER_66_216 VDD VSS sg13g2_decap_8
XFILLER_82_709 VDD VSS sg13g2_decap_8
XFILLER_86_84 VDD VSS sg13g2_decap_8
XFILLER_13_7 VDD VSS sg13g2_decap_8
XFILLER_62_400 VDD VSS sg13g2_decap_8
XFILLER_19_154 VDD VSS sg13g2_decap_8
XFILLER_90_731 VDD VSS sg13g2_decap_8
XFILLER_74_293 VDD VSS sg13g2_decap_8
XFILLER_63_956 VDD VSS sg13g2_decap_8
XFILLER_35_658 VDD VSS sg13g2_decap_8
XFILLER_16_861 VDD VSS sg13g2_decap_8
XFILLER_76_1060 VDD VSS sg13g2_fill_1
XFILLER_37_1022 VDD VSS sg13g2_decap_8
XFILLER_62_477 VDD VSS sg13g2_decap_8
XFILLER_15_371 VDD VSS sg13g2_decap_8
XFILLER_22_308 VDD VSS sg13g2_decap_8
XFILLER_34_168 VDD VSS sg13g2_decap_8
X_1902_ _1903_/A _1903_/B _1911_/A VDD VSS sg13g2_nor2_1
XFILLER_31_875 VDD VSS sg13g2_decap_8
X_1833_ _2248_/Q _2207_/Q _1850_/B VDD VSS sg13g2_nor2b_1
XFILLER_30_385 VDD VSS sg13g2_decap_8
X_1764_ _1940_/A _2227_/Q _2235_/Q VDD VSS sg13g2_xnor2_1
Xhold526 _2369_/Q VDD VSS hold526/X sg13g2_dlygate4sd3_1
Xhold515 _1711_/Y VDD VSS _1712_/B sg13g2_dlygate4sd3_1
Xhold504 _1695_/Y VDD VSS _1696_/B sg13g2_dlygate4sd3_1
XFILLER_7_581 VDD VSS sg13g2_decap_8
XFILLER_104_619 VDD VSS sg13g2_decap_8
Xhold537 _2203_/Q VDD VSS hold537/X sg13g2_dlygate4sd3_1
Xhold559 _2320_/Q VDD VSS hold559/X sg13g2_dlygate4sd3_1
X_1695_ _1694_/Y VDD _1695_/Y VSS _1724_/S hold503/X sg13g2_o21ai_1
Xhold548 _1614_/Y VDD VSS _1615_/B sg13g2_dlygate4sd3_1
XFILLER_83_1031 VDD VSS sg13g2_decap_8
XFILLER_98_820 VDD VSS sg13g2_decap_8
XFILLER_112_630 VDD VSS sg13g2_decap_8
XFILLER_97_352 VDD VSS sg13g2_fill_1
XFILLER_106_28 VDD VSS sg13g2_decap_8
XFILLER_44_1026 VDD VSS sg13g2_decap_8
X_2316_ _2316_/RESET_B VSS VDD _2316_/D _2316_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_85_503 VDD VSS sg13g2_decap_8
XFILLER_111_140 VDD VSS sg13g2_decap_8
XFILLER_39_920 VDD VSS sg13g2_decap_8
XFILLER_58_728 VDD VSS sg13g2_decap_8
XFILLER_100_847 VDD VSS sg13g2_decap_8
XFILLER_85_547 VDD VSS sg13g2_decap_8
X_2247_ _2247_/RESET_B VSS VDD _2247_/D _2247_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_997 VDD VSS sg13g2_decap_8
XFILLER_66_761 VDD VSS sg13g2_decap_8
XFILLER_38_474 VDD VSS sg13g2_decap_8
X_2178_ _2178_/RESET_B VSS VDD _2178_/D _2178_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_54_934 VDD VSS sg13g2_decap_8
XFILLER_80_241 VDD VSS sg13g2_decap_8
XFILLER_26_658 VDD VSS sg13g2_decap_8
XFILLER_15_14 VDD VSS sg13g2_decap_8
XFILLER_81_797 VDD VSS sg13g2_fill_2
XFILLER_53_477 VDD VSS sg13g2_decap_8
XFILLER_13_308 VDD VSS sg13g2_decap_8
XFILLER_40_105 VDD VSS sg13g2_decap_8
XFILLER_25_168 VDD VSS sg13g2_decap_8
XFILLER_90_1057 VDD VSS sg13g2_decap_4
X_2173__194 VDD VSS _2173_/RESET_B sg13g2_tiehi
XFILLER_22_875 VDD VSS sg13g2_decap_8
XFILLER_31_35 VDD VSS sg13g2_decap_8
XFILLER_21_385 VDD VSS sg13g2_decap_8
XFILLER_107_402 VDD VSS sg13g2_decap_8
XFILLER_5_518 VDD VSS sg13g2_decap_8
XFILLER_108_969 VDD VSS sg13g2_decap_8
XFILLER_107_479 VDD VSS sg13g2_decap_4
XFILLER_1_735 VDD VSS sg13g2_decap_8
Xout_data_pads\[0\].out_data_pad _2366_/Q IOVDD IOVSS out_data_PADs[0] VDD VSS sg13g2_IOPadOut30mA
XFILLER_103_630 VDD VSS sg13g2_decap_8
XFILLER_0_245 VDD VSS sg13g2_decap_8
XFILLER_88_363 VDD VSS sg13g2_fill_1
XFILLER_102_140 VDD VSS sg13g2_decap_8
XFILLER_49_739 VDD VSS sg13g2_decap_8
XFILLER_102_184 VDD VSS sg13g2_fill_1
XFILLER_56_32 VDD VSS sg13g2_fill_1
XFILLER_56_21 VDD VSS sg13g2_decap_8
XFILLER_99_1060 VDD VSS sg13g2_fill_1
XFILLER_91_528 VDD VSS sg13g2_decap_8
XFILLER_57_772 VDD VSS sg13g2_decap_8
XFILLER_29_441 VDD VSS sg13g2_decap_8
XFILLER_56_76 VDD VSS sg13g2_decap_8
XFILLER_45_989 VDD VSS sg13g2_decap_8
XFILLER_17_658 VDD VSS sg13g2_decap_8
XFILLER_71_263 VDD VSS sg13g2_fill_2
XFILLER_72_42 VDD VSS sg13g2_decap_8
XFILLER_16_168 VDD VSS sg13g2_decap_8
XFILLER_31_105 VDD VSS sg13g2_decap_8
XFILLER_44_488 VDD VSS sg13g2_decap_8
XFILLER_8_301 VDD VSS sg13g2_decap_8
XFILLER_13_875 VDD VSS sg13g2_decap_8
XFILLER_40_683 VDD VSS sg13g2_decap_8
XFILLER_12_385 VDD VSS sg13g2_decap_8
XFILLER_9_868 VDD VSS sg13g2_decap_8
XFILLER_8_378 VDD VSS sg13g2_decap_8
XFILLER_99_639 VDD VSS sg13g2_decap_8
XFILLER_98_105 VDD VSS sg13g2_decap_8
XFILLER_4_595 VDD VSS sg13g2_decap_8
X_1480_ _1602_/B VDD _1480_/Y VSS _1388_/A _1481_/A2 sg13g2_o21ai_1
XFILLER_95_801 VDD VSS sg13g2_decap_8
XFILLER_79_341 VDD VSS sg13g2_decap_8
XFILLER_79_363 VDD VSS sg13g2_decap_8
XFILLER_67_525 VDD VSS sg13g2_decap_8
XFILLER_39_238 VDD VSS sg13g2_decap_8
X_2101_ _2101_/A _2101_/B _2352_/D VDD VSS sg13g2_nor2_1
XFILLER_95_889 VDD VSS sg13g2_decap_8
X_2032_ _2071_/B _2156_/A _2082_/B VDD VSS sg13g2_nor2_1
XFILLER_94_377 VDD VSS sg13g2_decap_8
XFILLER_82_506 VDD VSS sg13g2_decap_8
XFILLER_48_761 VDD VSS sg13g2_decap_8
XFILLER_36_945 VDD VSS sg13g2_decap_8
XFILLER_47_271 VDD VSS sg13g2_decap_8
XFILLER_51_904 VDD VSS sg13g2_decap_8
XFILLER_35_455 VDD VSS sg13g2_decap_8
XFILLER_63_786 VDD VSS sg13g2_decap_8
XFILLER_22_105 VDD VSS sg13g2_decap_8
XFILLER_90_594 VDD VSS sg13g2_decap_8
XFILLER_50_458 VDD VSS sg13g2_decap_8
XFILLER_87_0 VDD VSS sg13g2_decap_8
XFILLER_31_672 VDD VSS sg13g2_decap_8
XFILLER_30_182 VDD VSS sg13g2_decap_8
X_1816_ _1901_/A _1930_/A _1816_/B VDD VSS sg13g2_nand2_1
XFILLER_50_1052 VDD VSS sg13g2_decap_8
XFILLER_7_70 VDD VSS sg13g2_decap_8
XFILLER_11_1036 VDD VSS sg13g2_decap_8
Xhold301 _2358_/Q VDD VSS _1502_/A sg13g2_dlygate4sd3_1
XFILLER_105_917 VDD VSS sg13g2_decap_8
Xhold323 _1274_/Y VDD VSS _1275_/A sg13g2_dlygate4sd3_1
Xhold312 _2170_/Q VDD VSS hold312/X sg13g2_dlygate4sd3_1
Xhold334 _2181_/Q VDD VSS hold334/X sg13g2_dlygate4sd3_1
XFILLER_104_405 VDD VSS sg13g2_fill_1
X_1747_ _2240_/Q _2232_/Q _1749_/A VDD VSS sg13g2_nor2b_1
Xhold345 _2166_/Q VDD VSS hold345/X sg13g2_dlygate4sd3_1
Xhold367 _1340_/Y VDD VSS _1341_/A sg13g2_dlygate4sd3_1
Xhold356 _1288_/Y VDD VSS _1289_/A sg13g2_dlygate4sd3_1
Xhold378 _1318_/Y VDD VSS _1319_/A sg13g2_dlygate4sd3_1
XFILLER_89_105 VDD VSS sg13g2_decap_8
X_1678_ _1681_/A _1678_/B _1679_/B VDD VSS sg13g2_nor2_1
Xhold389 _2188_/Q VDD VSS hold389/X sg13g2_dlygate4sd3_1
XFILLER_86_823 VDD VSS sg13g2_decap_8
XFILLER_58_525 VDD VSS sg13g2_decap_8
XFILLER_100_644 VDD VSS sg13g2_decap_8
XFILLER_97_193 VDD VSS sg13g2_decap_8
XFILLER_85_355 VDD VSS sg13g2_decap_8
XFILLER_73_517 VDD VSS sg13g2_decap_8
XFILLER_27_945 VDD VSS sg13g2_decap_8
XFILLER_66_580 VDD VSS sg13g2_fill_2
XFILLER_39_794 VDD VSS sg13g2_decap_8
XFILLER_26_35 VDD VSS sg13g2_decap_8
XFILLER_26_455 VDD VSS sg13g2_decap_8
XFILLER_53_252 VDD VSS sg13g2_fill_2
XFILLER_13_105 VDD VSS sg13g2_decap_8
XFILLER_81_594 VDD VSS sg13g2_decap_8
XFILLER_42_959 VDD VSS sg13g2_decap_8
XFILLER_53_285 VDD VSS sg13g2_decap_8
XFILLER_41_458 VDD VSS sg13g2_decap_8
XFILLER_107_1031 VDD VSS sg13g2_decap_8
XFILLER_10_812 VDD VSS sg13g2_decap_8
XFILLER_50_981 VDD VSS sg13g2_decap_8
XFILLER_22_672 VDD VSS sg13g2_decap_8
XFILLER_42_56 VDD VSS sg13g2_decap_8
XFILLER_6_805 VDD VSS sg13g2_decap_8
XFILLER_21_182 VDD VSS sg13g2_decap_8
XFILLER_5_315 VDD VSS sg13g2_decap_8
XFILLER_10_889 VDD VSS sg13g2_decap_8
XFILLER_108_766 VDD VSS sg13g2_decap_8
XFILLER_107_298 VDD VSS sg13g2_decap_8
XFILLER_104_950 VDD VSS sg13g2_decap_8
XFILLER_1_532 VDD VSS sg13g2_decap_8
XFILLER_3_28 VDD VSS sg13g2_decap_8
XFILLER_77_823 VDD VSS sg13g2_decap_8
XFILLER_95_119 VDD VSS sg13g2_decap_8
XFILLER_27_1043 VDD VSS sg13g2_decap_8
XFILLER_49_514 VDD VSS sg13g2_decap_8
XFILLER_77_856 VDD VSS sg13g2_decap_8
XFILLER_103_482 VDD VSS sg13g2_decap_8
XFILLER_49_558 VDD VSS sg13g2_decap_8
XFILLER_67_42 VDD VSS sg13g2_decap_8
XFILLER_49_525 VDD VSS sg13g2_fill_1
XFILLER_92_826 VDD VSS sg13g2_decap_8
XFILLER_18_945 VDD VSS sg13g2_decap_8
XFILLER_72_550 VDD VSS sg13g2_decap_8
XFILLER_17_455 VDD VSS sg13g2_decap_8
XFILLER_83_63 VDD VSS sg13g2_decap_8
XFILLER_44_252 VDD VSS sg13g2_fill_1
XFILLER_73_1030 VDD VSS sg13g2_decap_8
XFILLER_33_959 VDD VSS sg13g2_decap_8
XFILLER_60_778 VDD VSS sg13g2_decap_8
XFILLER_20_609 VDD VSS sg13g2_decap_8
XFILLER_32_469 VDD VSS sg13g2_decap_8
XFILLER_80_7 VDD VSS sg13g2_decap_8
XFILLER_34_1036 VDD VSS sg13g2_decap_8
XFILLER_13_672 VDD VSS sg13g2_decap_8
XFILLER_12_182 VDD VSS sg13g2_decap_8
XFILLER_9_665 VDD VSS sg13g2_decap_8
XFILLER_40_491 VDD VSS sg13g2_decap_8
XFILLER_8_175 VDD VSS sg13g2_decap_8
X_1601_ _1601_/Y _1638_/S _1607_/A VDD VSS sg13g2_nand2_1
X_1532_ _1531_/Y VDD _1532_/Y VSS _1592_/A _1529_/Y sg13g2_o21ai_1
XFILLER_5_882 VDD VSS sg13g2_decap_8
XFILLER_102_909 VDD VSS sg13g2_decap_8
XFILLER_87_609 VDD VSS sg13g2_decap_8
XFILLER_99_469 VDD VSS sg13g2_decap_8
X_1463_ _1463_/A _1463_/B _1463_/Y VDD VSS sg13g2_nor2_1
XFILLER_4_392 VDD VSS sg13g2_decap_8
XFILLER_80_1001 VDD VSS sg13g2_decap_8
XFILLER_110_942 VDD VSS sg13g2_decap_8
X_1394_ VDD _2219_/D _1394_/A VSS sg13g2_inv_1
XFILLER_41_1007 VDD VSS sg13g2_decap_8
XFILLER_68_834 VDD VSS sg13g2_decap_8
XFILLER_67_322 VDD VSS sg13g2_decap_8
XFILLER_83_815 VDD VSS sg13g2_decap_8
XFILLER_95_686 VDD VSS sg13g2_decap_8
X_2015_ _2015_/Y _2022_/S _2015_/B VDD VSS sg13g2_nand2_1
XFILLER_94_196 VDD VSS sg13g2_decap_8
XFILLER_36_742 VDD VSS sg13g2_decap_8
X_2239__264 VDD VSS _2239_/RESET_B sg13g2_tiehi
XFILLER_35_252 VDD VSS sg13g2_decap_8
XFILLER_24_959 VDD VSS sg13g2_decap_8
XFILLER_11_609 VDD VSS sg13g2_decap_8
XFILLER_23_469 VDD VSS sg13g2_decap_8
XFILLER_10_119 VDD VSS sg13g2_decap_8
XFILLER_3_819 VDD VSS sg13g2_decap_8
XFILLER_105_714 VDD VSS sg13g2_decap_8
XFILLER_104_202 VDD VSS sg13g2_decap_8
XFILLER_2_329 VDD VSS sg13g2_decap_8
XFILLER_104_224 VDD VSS sg13g2_decap_8
XFILLER_77_119 VDD VSS sg13g2_decap_8
XFILLER_101_942 VDD VSS sg13g2_decap_8
XFILLER_58_344 VDD VSS sg13g2_decap_8
XFILLER_86_686 VDD VSS sg13g2_decap_8
XFILLER_100_496 VDD VSS sg13g2_decap_8
XFILLER_85_185 VDD VSS sg13g2_decap_8
XFILLER_58_399 VDD VSS sg13g2_decap_8
XFILLER_2_1001 VDD VSS sg13g2_decap_8
XFILLER_37_56 VDD VSS sg13g2_decap_8
XFILLER_46_517 VDD VSS sg13g2_decap_8
XFILLER_73_358 VDD VSS sg13g2_decap_8
XFILLER_39_591 VDD VSS sg13g2_decap_8
XFILLER_27_742 VDD VSS sg13g2_decap_8
XFILLER_61_509 VDD VSS sg13g2_fill_2
XFILLER_26_252 VDD VSS sg13g2_decap_8
XFILLER_42_756 VDD VSS sg13g2_decap_8
XFILLER_15_959 VDD VSS sg13g2_decap_8
XFILLER_14_469 VDD VSS sg13g2_decap_8
XFILLER_53_55 VDD VSS sg13g2_decap_8
XFILLER_41_255 VDD VSS sg13g2_decap_8
XFILLER_6_602 VDD VSS sg13g2_decap_8
XFILLER_5_112 VDD VSS sg13g2_decap_8
XFILLER_10_686 VDD VSS sg13g2_decap_8
XFILLER_6_679 VDD VSS sg13g2_decap_8
XFILLER_108_563 VDD VSS sg13g2_decap_8
XFILLER_5_189 VDD VSS sg13g2_decap_8
XFILLER_64_1007 VDD VSS sg13g2_fill_2
XFILLER_111_728 VDD VSS sg13g2_decap_8
XFILLER_96_406 VDD VSS sg13g2_decap_8
XFILLER_78_63 VDD VSS sg13g2_decap_8
XFILLER_110_238 VDD VSS sg13g2_decap_8
XFILLER_2_896 VDD VSS sg13g2_decap_8
XFILLER_77_653 VDD VSS sg13g2_decap_8
XFILLER_49_344 VDD VSS sg13g2_decap_8
XFILLER_40_1040 VDD VSS sg13g2_decap_8
XFILLER_64_314 VDD VSS sg13g2_decap_8
XFILLER_37_539 VDD VSS sg13g2_decap_8
XFILLER_76_196 VDD VSS sg13g2_decap_8
XFILLER_94_84 VDD VSS sg13g2_decap_8
XFILLER_18_742 VDD VSS sg13g2_decap_8
XFILLER_92_689 VDD VSS sg13g2_decap_8
XFILLER_17_252 VDD VSS sg13g2_decap_8
XFILLER_91_199 VDD VSS sg13g2_decap_8
XFILLER_72_391 VDD VSS sg13g2_fill_1
XFILLER_72_380 VDD VSS sg13g2_decap_8
XFILLER_33_756 VDD VSS sg13g2_decap_8
XFILLER_60_531 VDD VSS sg13g2_decap_8
XFILLER_20_406 VDD VSS sg13g2_decap_8
XFILLER_32_266 VDD VSS sg13g2_decap_8
XFILLER_9_462 VDD VSS sg13g2_decap_8
X_2345__123 VDD VSS _2345_/RESET_B sg13g2_tiehi
XFILLER_88_907 VDD VSS sg13g2_decap_8
X_1515_ _1260_/A VDD _1515_/Y VSS _1503_/X _1514_/Y sg13g2_o21ai_1
XFILLER_101_205 VDD VSS sg13g2_decap_4
XFILLER_96_940 VDD VSS sg13g2_decap_8
XFILLER_101_227 VDD VSS sg13g2_decap_8
X_1446_ VDD VSS _1265_/B _1228_/A _1218_/Y _1193_/Y _1446_/Y _1501_/A sg13g2_a221oi_1
X_1377_ _1377_/Y _1377_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_83_612 VDD VSS sg13g2_decap_8
XFILLER_95_494 VDD VSS sg13g2_fill_1
XFILLER_95_483 VDD VSS sg13g2_decap_8
XFILLER_67_174 VDD VSS sg13g2_decap_8
XFILLER_28_539 VDD VSS sg13g2_decap_8
XFILLER_83_656 VDD VSS sg13g2_fill_1
XFILLER_55_336 VDD VSS sg13g2_decap_8
XFILLER_70_306 VDD VSS sg13g2_decap_8
X_2356__274 VDD VSS _2356_/RESET_B sg13g2_tiehi
XFILLER_70_339 VDD VSS sg13g2_fill_2
XFILLER_63_380 VDD VSS sg13g2_decap_8
XFILLER_24_756 VDD VSS sg13g2_decap_8
XFILLER_11_406 VDD VSS sg13g2_decap_8
XFILLER_51_586 VDD VSS sg13g2_decap_8
XFILLER_23_14 VDD VSS sg13g2_decap_8
XFILLER_23_266 VDD VSS sg13g2_decap_8
XFILLER_104_1034 VDD VSS sg13g2_decap_8
XFILLER_20_973 VDD VSS sg13g2_decap_8
XFILLER_3_616 VDD VSS sg13g2_decap_8
X_2324__218 VDD VSS _2324_/RESET_B sg13g2_tiehi
XFILLER_105_533 VDD VSS sg13g2_decap_8
XFILLER_2_126 VDD VSS sg13g2_decap_8
XFILLER_79_929 VDD VSS sg13g2_fill_1
XFILLER_105_588 VDD VSS sg13g2_decap_8
XFILLER_78_417 VDD VSS sg13g2_decap_8
XFILLER_63_1051 VDD VSS sg13g2_decap_8
XFILLER_59_664 VDD VSS sg13g2_decap_8
XFILLER_101_772 VDD VSS sg13g2_decap_8
XFILLER_86_461 VDD VSS sg13g2_decap_8
XFILLER_24_1057 VDD VSS sg13g2_decap_4
XFILLER_19_539 VDD VSS sg13g2_decap_8
XFILLER_74_667 VDD VSS sg13g2_decap_8
XFILLER_100_282 VDD VSS sg13g2_decap_4
XFILLER_100_293 VDD VSS sg13g2_decap_8
XFILLER_47_859 VDD VSS sg13g2_decap_8
XFILLER_64_21 VDD VSS sg13g2_decap_8
XFILLER_46_347 VDD VSS sg13g2_fill_2
XFILLER_62_829 VDD VSS sg13g2_decap_8
XFILLER_55_881 VDD VSS sg13g2_decap_8
XFILLER_46_369 VDD VSS sg13g2_fill_1
XFILLER_54_380 VDD VSS sg13g2_decap_4
XFILLER_42_520 VDD VSS sg13g2_decap_4
XFILLER_42_564 VDD VSS sg13g2_fill_1
XFILLER_15_756 VDD VSS sg13g2_decap_8
XFILLER_70_1011 VDD VSS sg13g2_decap_8
XFILLER_80_42 VDD VSS sg13g2_decap_8
XFILLER_14_266 VDD VSS sg13g2_decap_8
XFILLER_9_49 VDD VSS sg13g2_decap_8
XFILLER_70_1044 VDD VSS sg13g2_decap_8
Xfanout70 _2106_/A _1228_/A VDD VSS sg13g2_buf_1
XFILLER_11_973 VDD VSS sg13g2_decap_8
XFILLER_109_861 VDD VSS sg13g2_decap_8
XFILLER_10_483 VDD VSS sg13g2_decap_8
XFILLER_13_91 VDD VSS sg13g2_decap_8
XFILLER_7_966 VDD VSS sg13g2_decap_8
XFILLER_108_360 VDD VSS sg13g2_decap_4
XFILLER_6_476 VDD VSS sg13g2_decap_8
XFILLER_89_84 VDD VSS sg13g2_decap_8
XFILLER_97_715 VDD VSS sg13g2_decap_8
XFILLER_96_203 VDD VSS sg13g2_decap_8
XFILLER_9_1029 VDD VSS sg13g2_decap_8
XFILLER_43_7 VDD VSS sg13g2_decap_8
XFILLER_97_737 VDD VSS sg13g2_decap_4
XFILLER_111_525 VDD VSS sg13g2_decap_8
X_1300_ _1300_/Y _1344_/B1 hold308/X _1344_/A2 _2344_/Q VDD VSS sg13g2_a22oi_1
XFILLER_2_693 VDD VSS sg13g2_decap_8
X_2280_ _2280_/RESET_B VSS VDD _2280_/D _2280_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_78_951 VDD VSS sg13g2_decap_8
X_1231_ _1234_/B _1365_/B _2355_/Q VDD VSS sg13g2_nand2_1
XFILLER_77_461 VDD VSS sg13g2_decap_8
XFILLER_93_965 VDD VSS sg13g2_decap_8
XFILLER_65_634 VDD VSS sg13g2_decap_8
XFILLER_65_645 VDD VSS sg13g2_fill_2
XFILLER_37_336 VDD VSS sg13g2_decap_8
XFILLER_49_196 VDD VSS sg13g2_decap_8
XFILLER_65_689 VDD VSS sg13g2_decap_8
XFILLER_80_637 VDD VSS sg13g2_decap_8
XFILLER_80_648 VDD VSS sg13g2_fill_1
XFILLER_64_199 VDD VSS sg13g2_fill_1
XFILLER_61_851 VDD VSS sg13g2_decap_8
XFILLER_33_553 VDD VSS sg13g2_decap_8
XFILLER_20_203 VDD VSS sg13g2_decap_8
X_1995_ _1995_/A _1995_/B _1995_/C _1995_/X VDD VSS sg13g2_or3_1
XFILLER_109_28 VDD VSS sg13g2_decap_8
XFILLER_106_319 VDD VSS sg13g2_decap_8
XFILLER_47_1013 VDD VSS sg13g2_decap_8
XFILLER_102_514 VDD VSS sg13g2_decap_8
XFILLER_87_269 VDD VSS sg13g2_decap_8
X_1429_ _1429_/A _1429_/B _1429_/Y VDD VSS sg13g2_nor2_1
XFILLER_69_995 VDD VSS sg13g2_fill_2
XFILLER_56_623 VDD VSS sg13g2_decap_8
XFILLER_29_826 VDD VSS sg13g2_decap_8
XFILLER_18_14 VDD VSS sg13g2_decap_8
XFILLER_84_954 VDD VSS sg13g2_decap_8
XFILLER_83_431 VDD VSS sg13g2_decap_8
XFILLER_68_494 VDD VSS sg13g2_decap_8
XFILLER_55_133 VDD VSS sg13g2_decap_8
XFILLER_28_336 VDD VSS sg13g2_decap_8
XFILLER_84_987 VDD VSS sg13g2_decap_8
XFILLER_71_626 VDD VSS sg13g2_decap_8
XFILLER_44_818 VDD VSS sg13g2_decap_8
XFILLER_43_306 VDD VSS sg13g2_fill_2
XIO_BOND_in_data_pads\[0\].in_data_pad in_data_PADs[0] bondpad_70x70
XFILLER_93_1011 VDD VSS sg13g2_decap_8
XFILLER_70_147 VDD VSS sg13g2_decap_8
XFILLER_24_553 VDD VSS sg13g2_decap_8
XFILLER_34_35 VDD VSS sg13g2_decap_8
XFILLER_11_203 VDD VSS sg13g2_decap_8
Xclkload1 clkload1/Y clkload1/A VDD VSS sg13g2_inv_2
XFILLER_20_770 VDD VSS sg13g2_decap_8
XFILLER_109_168 VDD VSS sg13g2_decap_8
XFILLER_30_1050 VDD VSS sg13g2_decap_8
XFILLER_4_903 VDD VSS sg13g2_decap_8
XFILLER_106_853 VDD VSS sg13g2_decap_8
XFILLER_3_413 VDD VSS sg13g2_decap_8
XFILLER_79_715 VDD VSS sg13g2_decap_8
XFILLER_105_330 VDD VSS sg13g2_decap_8
XFILLER_59_21 VDD VSS sg13g2_decap_8
X_2183__174 VDD VSS _2183_/RESET_B sg13g2_tiehi
XFILLER_47_623 VDD VSS sg13g2_decap_8
XFILLER_59_483 VDD VSS sg13g2_decap_8
XFILLER_59_450 VDD VSS sg13g2_decap_8
XFILLER_101_580 VDD VSS sg13g2_decap_8
XFILLER_74_431 VDD VSS sg13g2_decap_8
XFILLER_75_42 VDD VSS sg13g2_decap_8
XFILLER_19_336 VDD VSS sg13g2_decap_8
XFILLER_90_902 VDD VSS sg13g2_decap_8
XFILLER_74_475 VDD VSS sg13g2_decap_4
XFILLER_74_486 VDD VSS sg13g2_decap_8
XFILLER_62_648 VDD VSS sg13g2_decap_8
XFILLER_46_199 VDD VSS sg13g2_decap_8
XFILLER_15_553 VDD VSS sg13g2_decap_8
XFILLER_61_136 VDD VSS sg13g2_decap_8
XFILLER_91_63 VDD VSS sg13g2_decap_8
XFILLER_43_884 VDD VSS sg13g2_decap_8
XFILLER_42_350 VDD VSS sg13g2_decap_8
X_1780_ _1780_/Y _2220_/Q _2212_/Q VDD VSS sg13g2_nand2b_1
XFILLER_30_567 VDD VSS sg13g2_decap_8
XFILLER_11_770 VDD VSS sg13g2_decap_8
XFILLER_10_280 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_7_763 VDD VSS sg13g2_decap_8
XFILLER_6_273 VDD VSS sg13g2_decap_8
XFILLER_112_812 VDD VSS sg13g2_decap_8
X_2332_ _2332_/RESET_B VSS VDD _2332_/D _2332_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_69_225 VDD VSS sg13g2_fill_1
XFILLER_3_980 VDD VSS sg13g2_decap_8
XFILLER_97_556 VDD VSS sg13g2_decap_8
XFILLER_111_322 VDD VSS sg13g2_decap_8
XFILLER_2_490 VDD VSS sg13g2_decap_8
XFILLER_112_889 VDD VSS sg13g2_decap_8
XFILLER_66_921 VDD VSS sg13g2_decap_8
X_2263_ _2263_/RESET_B VSS VDD _2263_/D _2263_/Q clkload1/A sg13g2_dfrbpq_1
X_2194_ _2194_/RESET_B VSS VDD _2194_/D _2194_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_111_399 VDD VSS sg13g2_decap_8
XFILLER_77_280 VDD VSS sg13g2_decap_8
X_1214_ VDD _1214_/Y _2245_/Q VSS sg13g2_inv_1
XFILLER_37_133 VDD VSS sg13g2_decap_8
XFILLER_93_773 VDD VSS sg13g2_decap_8
X_2273__209 VDD VSS _2273_/RESET_B sg13g2_tiehi
XFILLER_38_667 VDD VSS sg13g2_decap_8
XFILLER_81_946 VDD VSS sg13g2_decap_8
XFILLER_77_1028 VDD VSS sg13g2_decap_8
XFILLER_80_467 VDD VSS sg13g2_decap_8
XFILLER_34_840 VDD VSS sg13g2_decap_8
XFILLER_61_670 VDD VSS sg13g2_fill_2
X_2353__288 VDD VSS _2353_/RESET_B sg13g2_tiehi
XFILLER_33_350 VDD VSS sg13g2_decap_8
XFILLER_21_567 VDD VSS sg13g2_decap_8
XFILLER_14_1001 VDD VSS sg13g2_decap_8
X_1978_ _1978_/A _1978_/B _1978_/C _1982_/C VDD VSS sg13g2_or3_1
XFILLER_101_1048 VDD VSS sg13g2_decap_8
XFILLER_106_105 VDD VSS sg13g2_decap_8
XFILLER_101_1059 VDD VSS sg13g2_fill_2
XFILLER_107_639 VDD VSS sg13g2_decap_8
XFILLER_1_917 VDD VSS sg13g2_decap_8
XFILLER_0_427 VDD VSS sg13g2_decap_8
XFILLER_103_856 VDD VSS sg13g2_fill_1
XFILLER_29_35 VDD VSS sg13g2_decap_8
XFILLER_48_409 VDD VSS sg13g2_decap_8
XFILLER_88_589 VDD VSS sg13g2_fill_1
XFILLER_60_1032 VDD VSS sg13g2_decap_8
XFILLER_84_740 VDD VSS sg13g2_decap_8
XFILLER_57_943 VDD VSS sg13g2_fill_1
XFILLER_29_623 VDD VSS sg13g2_decap_8
XFILLER_68_291 VDD VSS sg13g2_decap_8
XFILLER_90_209 VDD VSS sg13g2_decap_4
XFILLER_28_133 VDD VSS sg13g2_decap_8
XFILLER_56_497 VDD VSS sg13g2_decap_8
XFILLER_45_56 VDD VSS sg13g2_decap_8
XFILLER_71_467 VDD VSS sg13g2_decap_8
XFILLER_25_840 VDD VSS sg13g2_decap_8
XFILLER_43_147 VDD VSS sg13g2_decap_8
XFILLER_24_350 VDD VSS sg13g2_decap_8
XFILLER_101_84 VDD VSS sg13g2_decap_8
XFILLER_40_865 VDD VSS sg13g2_decap_8
XFILLER_12_567 VDD VSS sg13g2_decap_8
XFILLER_61_77 VDD VSS sg13g2_decap_4
XFILLER_61_99 VDD VSS sg13g2_fill_1
XFILLER_6_28 VDD VSS sg13g2_decap_8
XFILLER_4_700 VDD VSS sg13g2_decap_8
XFILLER_3_210 VDD VSS sg13g2_decap_8
XFILLER_106_650 VDD VSS sg13g2_decap_8
XFILLER_4_777 VDD VSS sg13g2_decap_8
XFILLER_79_512 VDD VSS sg13g2_decap_8
XFILLER_112_119 VDD VSS sg13g2_decap_8
XFILLER_3_287 VDD VSS sg13g2_decap_8
XFILLER_10_70 VDD VSS sg13g2_decap_8
XFILLER_67_707 VDD VSS sg13g2_fill_1
XFILLER_94_515 VDD VSS sg13g2_decap_8
XFILLER_86_63 VDD VSS sg13g2_decap_8
XFILLER_59_291 VDD VSS sg13g2_decap_8
XFILLER_0_994 VDD VSS sg13g2_decap_8
XFILLER_63_902 VDD VSS sg13g2_decap_8
XFILLER_19_133 VDD VSS sg13g2_decap_8
XFILLER_47_442 VDD VSS sg13g2_fill_2
XFILLER_90_710 VDD VSS sg13g2_decap_8
XFILLER_74_272 VDD VSS sg13g2_decap_8
XFILLER_35_637 VDD VSS sg13g2_decap_8
XFILLER_37_1001 VDD VSS sg13g2_decap_8
XFILLER_62_456 VDD VSS sg13g2_decap_8
XFILLER_16_840 VDD VSS sg13g2_decap_8
XFILLER_34_147 VDD VSS sg13g2_decap_8
XFILLER_90_787 VDD VSS sg13g2_decap_8
XFILLER_50_618 VDD VSS sg13g2_fill_1
XFILLER_43_681 VDD VSS sg13g2_decap_8
XFILLER_15_350 VDD VSS sg13g2_decap_8
X_1901_ _1901_/B _1901_/A _1903_/B VDD VSS sg13g2_xor2_1
XFILLER_31_854 VDD VSS sg13g2_decap_8
XFILLER_42_191 VDD VSS sg13g2_decap_8
X_1832_ _1852_/B _2249_/Q _2208_/Q VDD VSS sg13g2_nand2b_1
XFILLER_30_364 VDD VSS sg13g2_decap_8
X_1763_ _1948_/A _1763_/A _1763_/B VDD VSS sg13g2_xnor2_1
XFILLER_7_560 VDD VSS sg13g2_decap_8
Xhold516 _1712_/Y VDD VSS _2317_/D sg13g2_dlygate4sd3_1
X_1694_ _1694_/Y _1724_/S _1698_/A VDD VSS sg13g2_nand2_1
Xhold505 _1696_/Y VDD VSS _2314_/D sg13g2_dlygate4sd3_1
Xhold527 _2290_/Q VDD VSS hold527/X sg13g2_dlygate4sd3_1
Xhold538 _2371_/Q VDD VSS hold538/X sg13g2_dlygate4sd3_1
Xhold549 _1615_/Y VDD VSS _2292_/D sg13g2_dlygate4sd3_1
XFILLER_103_119 VDD VSS sg13g2_decap_8
XFILLER_44_1005 VDD VSS sg13g2_decap_8
XFILLER_58_707 VDD VSS sg13g2_decap_8
XFILLER_32_0 VDD VSS sg13g2_decap_8
X_2315_ _2315_/RESET_B VSS VDD _2315_/D _2315_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_112_686 VDD VSS sg13g2_decap_8
XFILLER_100_804 VDD VSS sg13g2_fill_2
XFILLER_98_898 VDD VSS sg13g2_decap_8
XFILLER_97_386 VDD VSS sg13g2_decap_8
XFILLER_85_526 VDD VSS sg13g2_decap_8
XFILLER_111_196 VDD VSS sg13g2_decap_8
X_2246_ _2246_/RESET_B VSS VDD _2246_/D _2246_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_57_239 VDD VSS sg13g2_decap_8
XFILLER_39_976 VDD VSS sg13g2_decap_8
XFILLER_54_913 VDD VSS sg13g2_decap_4
XFILLER_38_453 VDD VSS sg13g2_decap_8
X_2177_ _2177_/RESET_B VSS VDD _2177_/D _2177_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_66_784 VDD VSS sg13g2_fill_1
XFILLER_26_637 VDD VSS sg13g2_decap_8
XFILLER_81_743 VDD VSS sg13g2_decap_8
XFILLER_81_754 VDD VSS sg13g2_fill_2
XFILLER_80_220 VDD VSS sg13g2_decap_8
XFILLER_53_456 VDD VSS sg13g2_decap_8
XFILLER_25_147 VDD VSS sg13g2_decap_8
XFILLER_41_629 VDD VSS sg13g2_decap_8
XFILLER_90_1036 VDD VSS sg13g2_decap_8
XFILLER_22_854 VDD VSS sg13g2_decap_8
XFILLER_21_364 VDD VSS sg13g2_decap_8
XFILLER_31_14 VDD VSS sg13g2_decap_8
XFILLER_108_948 VDD VSS sg13g2_decap_8
XFILLER_110_7 VDD VSS sg13g2_decap_8
XFILLER_107_458 VDD VSS sg13g2_decap_8
XFILLER_1_714 VDD VSS sg13g2_decap_8
XFILLER_0_224 VDD VSS sg13g2_decap_8
XFILLER_89_887 VDD VSS sg13g2_decap_8
XFILLER_88_353 VDD VSS sg13g2_decap_4
XFILLER_76_526 VDD VSS sg13g2_decap_8
XFILLER_49_718 VDD VSS sg13g2_decap_8
XFILLER_29_420 VDD VSS sg13g2_decap_8
XFILLER_91_507 VDD VSS sg13g2_decap_8
XFILLER_57_751 VDD VSS sg13g2_decap_8
XFILLER_5_1043 VDD VSS sg13g2_decap_8
XFILLER_56_44 VDD VSS sg13g2_decap_8
XFILLER_84_592 VDD VSS sg13g2_decap_8
XFILLER_84_570 VDD VSS sg13g2_decap_4
XFILLER_17_637 VDD VSS sg13g2_decap_8
XFILLER_29_497 VDD VSS sg13g2_decap_8
XFILLER_72_754 VDD VSS sg13g2_fill_2
XFILLER_45_968 VDD VSS sg13g2_decap_8
XFILLER_16_147 VDD VSS sg13g2_decap_8
XFILLER_72_787 VDD VSS sg13g2_decap_8
XFILLER_72_21 VDD VSS sg13g2_decap_8
XFILLER_60_949 VDD VSS sg13g2_decap_8
XFILLER_44_467 VDD VSS sg13g2_decap_8
XFILLER_53_990 VDD VSS sg13g2_decap_8
XFILLER_13_854 VDD VSS sg13g2_decap_8
XFILLER_40_662 VDD VSS sg13g2_decap_8
XFILLER_12_364 VDD VSS sg13g2_decap_8
XFILLER_9_847 VDD VSS sg13g2_decap_8
XFILLER_8_357 VDD VSS sg13g2_decap_8
XFILLER_99_618 VDD VSS sg13g2_decap_8
XFILLER_21_91 VDD VSS sg13g2_decap_8
XFILLER_4_574 VDD VSS sg13g2_decap_8
XFILLER_79_320 VDD VSS sg13g2_decap_8
XFILLER_97_84 VDD VSS sg13g2_decap_8
XFILLER_67_504 VDD VSS sg13g2_decap_8
XFILLER_0_791 VDD VSS sg13g2_decap_8
XFILLER_39_217 VDD VSS sg13g2_decap_8
X_2100_ _2101_/B _2099_/X _2102_/B _2095_/A _2099_/A VDD VSS sg13g2_a22oi_1
X_2031_ _2031_/A _2089_/S _2031_/Y VDD VSS sg13g2_nor2b_1
XFILLER_94_367 VDD VSS sg13g2_fill_1
XFILLER_75_581 VDD VSS sg13g2_decap_8
XFILLER_36_924 VDD VSS sg13g2_decap_8
XFILLER_47_250 VDD VSS sg13g2_decap_8
XFILLER_63_765 VDD VSS sg13g2_decap_8
XFILLER_35_434 VDD VSS sg13g2_decap_8
XFILLER_50_437 VDD VSS sg13g2_decap_8
XFILLER_31_651 VDD VSS sg13g2_decap_8
XFILLER_30_161 VDD VSS sg13g2_decap_8
X_1815_ _1816_/B _1929_/B _1939_/B VDD VSS sg13g2_nand2_1
Xhold302 _2168_/Q VDD VSS hold302/X sg13g2_dlygate4sd3_1
X_1746_ VDD _1756_/B _1763_/B VSS sg13g2_inv_1
XFILLER_11_1015 VDD VSS sg13g2_decap_8
Xhold313 _1280_/Y VDD VSS _1281_/A sg13g2_dlygate4sd3_1
Xhold335 _1302_/Y VDD VSS _1303_/A sg13g2_dlygate4sd3_1
Xhold324 _2258_/Q VDD VSS _1195_/A sg13g2_dlygate4sd3_1
Xhold346 _1272_/Y VDD VSS _1273_/A sg13g2_dlygate4sd3_1
Xhold357 _2176_/Q VDD VSS hold357/X sg13g2_dlygate4sd3_1
Xhold368 _2198_/Q VDD VSS hold368/X sg13g2_dlygate4sd3_1
X_1677_ _1677_/A _1677_/B _1678_/B VDD VSS sg13g2_nor2_1
XFILLER_98_640 VDD VSS sg13g2_fill_2
Xhold379 _2163_/Q VDD VSS hold379/X sg13g2_dlygate4sd3_1
XFILLER_98_684 VDD VSS sg13g2_decap_8
XFILLER_86_802 VDD VSS sg13g2_decap_8
XFILLER_58_504 VDD VSS sg13g2_decap_8
XFILLER_100_623 VDD VSS sg13g2_decap_8
XFILLER_112_483 VDD VSS sg13g2_decap_8
XFILLER_97_172 VDD VSS sg13g2_decap_8
XFILLER_85_334 VDD VSS sg13g2_decap_8
XFILLER_100_689 VDD VSS sg13g2_decap_8
X_2229_ _2229__82/L_HI VSS VDD _2229_/D _2229_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_27_924 VDD VSS sg13g2_decap_8
XFILLER_39_773 VDD VSS sg13g2_decap_8
XFILLER_26_14 VDD VSS sg13g2_decap_8
XFILLER_66_592 VDD VSS sg13g2_decap_8
XFILLER_54_765 VDD VSS sg13g2_decap_8
XFILLER_26_434 VDD VSS sg13g2_decap_8
XFILLER_38_294 VDD VSS sg13g2_fill_1
XFILLER_81_573 VDD VSS sg13g2_decap_8
XFILLER_42_938 VDD VSS sg13g2_decap_8
XFILLER_54_787 VDD VSS sg13g2_fill_1
XFILLER_41_437 VDD VSS sg13g2_decap_8
XFILLER_107_1010 VDD VSS sg13g2_decap_8
XFILLER_50_960 VDD VSS sg13g2_decap_8
XFILLER_22_651 VDD VSS sg13g2_decap_8
XFILLER_42_35 VDD VSS sg13g2_decap_8
XFILLER_21_161 VDD VSS sg13g2_decap_8
XFILLER_10_868 VDD VSS sg13g2_decap_8
XFILLER_108_745 VDD VSS sg13g2_decap_8
XFILLER_107_266 VDD VSS sg13g2_decap_8
XFILLER_1_511 VDD VSS sg13g2_decap_8
XFILLER_66_1060 VDD VSS sg13g2_fill_1
XFILLER_77_802 VDD VSS sg13g2_decap_8
XFILLER_27_1022 VDD VSS sg13g2_decap_8
XFILLER_67_21 VDD VSS sg13g2_decap_8
XFILLER_88_161 VDD VSS sg13g2_decap_8
XFILLER_1_588 VDD VSS sg13g2_decap_8
XFILLER_49_537 VDD VSS sg13g2_decap_8
XFILLER_92_805 VDD VSS sg13g2_decap_8
XFILLER_67_98 VDD VSS sg13g2_decap_8
XFILLER_57_581 VDD VSS sg13g2_decap_8
XFILLER_64_529 VDD VSS sg13g2_decap_8
XFILLER_18_924 VDD VSS sg13g2_decap_8
XFILLER_91_348 VDD VSS sg13g2_decap_8
XFILLER_83_42 VDD VSS sg13g2_decap_8
XFILLER_17_434 VDD VSS sg13g2_decap_8
XFILLER_29_294 VDD VSS sg13g2_decap_8
XFILLER_33_938 VDD VSS sg13g2_decap_8
XFILLER_45_765 VDD VSS sg13g2_decap_8
XFILLER_45_776 VDD VSS sg13g2_fill_2
XFILLER_72_584 VDD VSS sg13g2_decap_8
XFILLER_32_448 VDD VSS sg13g2_decap_8
XFILLER_34_1015 VDD VSS sg13g2_decap_8
XFILLER_16_91 VDD VSS sg13g2_decap_8
XFILLER_13_651 VDD VSS sg13g2_decap_8
XFILLER_41_993 VDD VSS sg13g2_decap_8
XFILLER_12_161 VDD VSS sg13g2_decap_8
XFILLER_9_644 VDD VSS sg13g2_decap_8
XFILLER_73_7 VDD VSS sg13g2_decap_8
XFILLER_8_154 VDD VSS sg13g2_decap_8
X_1600_ _1607_/A _1637_/A _1600_/B VDD VSS sg13g2_xnor2_1
XFILLER_99_415 VDD VSS sg13g2_decap_4
XFILLER_99_404 VDD VSS sg13g2_fill_2
X_1531_ _1530_/Y VDD _1531_/Y VSS _1556_/S0 _2203_/Q sg13g2_o21ai_1
XFILLER_5_861 VDD VSS sg13g2_decap_8
XFILLER_99_448 VDD VSS sg13g2_decap_8
X_1462_ VSS VDD _1385_/Y _1463_/B _2250_/D _1461_/Y sg13g2_a21oi_1
XFILLER_4_371 VDD VSS sg13g2_decap_8
XFILLER_110_921 VDD VSS sg13g2_decap_8
XFILLER_80_1057 VDD VSS sg13g2_decap_4
XFILLER_95_610 VDD VSS sg13g2_decap_4
X_1393_ _1394_/A _1392_/Y hold550/X _1392_/B _1364_/A VDD VSS sg13g2_a22oi_1
XFILLER_79_161 VDD VSS sg13g2_decap_4
X_2308__81 VDD VSS _2308__81/L_HI sg13g2_tiehi
XFILLER_67_301 VDD VSS sg13g2_decap_8
XFILLER_95_665 VDD VSS sg13g2_decap_8
XFILLER_110_998 VDD VSS sg13g2_decap_8
XFILLER_82_315 VDD VSS sg13g2_fill_1
XFILLER_36_721 VDD VSS sg13g2_decap_8
XFILLER_55_529 VDD VSS sg13g2_decap_8
X_2014_ _2022_/S _2015_/B _2014_/X VDD VSS sg13g2_and2_1
XFILLER_35_231 VDD VSS sg13g2_decap_8
XFILLER_91_882 VDD VSS sg13g2_fill_2
XFILLER_24_938 VDD VSS sg13g2_decap_8
XFILLER_63_573 VDD VSS sg13g2_decap_8
XFILLER_36_798 VDD VSS sg13g2_decap_8
XFILLER_63_584 VDD VSS sg13g2_decap_4
XFILLER_23_448 VDD VSS sg13g2_decap_8
XFILLER_50_223 VDD VSS sg13g2_fill_2
XFILLER_51_779 VDD VSS sg13g2_decap_8
XFILLER_50_245 VDD VSS sg13g2_decap_8
XFILLER_12_49 VDD VSS sg13g2_decap_8
X_1729_ _2229_/Q _2237_/Q _1729_/Y VDD VSS sg13g2_nor2b_1
XFILLER_2_308 VDD VSS sg13g2_decap_8
XFILLER_101_921 VDD VSS sg13g2_fill_1
XFILLER_99_993 VDD VSS sg13g2_decap_8
XFILLER_59_857 VDD VSS sg13g2_decap_8
XFILLER_59_824 VDD VSS sg13g2_fill_2
XFILLER_58_323 VDD VSS sg13g2_decap_8
XFILLER_86_665 VDD VSS sg13g2_decap_8
XFILLER_112_280 VDD VSS sg13g2_decap_8
XFILLER_74_849 VDD VSS sg13g2_decap_4
XFILLER_100_475 VDD VSS sg13g2_fill_1
XFILLER_85_164 VDD VSS sg13g2_decap_8
XFILLER_39_570 VDD VSS sg13g2_decap_8
XFILLER_27_721 VDD VSS sg13g2_decap_8
XFILLER_37_35 VDD VSS sg13g2_decap_8
XFILLER_73_337 VDD VSS sg13g2_decap_8
XFILLER_26_231 VDD VSS sg13g2_decap_8
XFILLER_96_1053 VDD VSS sg13g2_decap_8
XFILLER_57_1004 VDD VSS sg13g2_fill_2
XFILLER_54_573 VDD VSS sg13g2_decap_4
XFILLER_2_1057 VDD VSS sg13g2_decap_4
XFILLER_82_893 VDD VSS sg13g2_decap_8
XFILLER_81_370 VDD VSS sg13g2_fill_1
XFILLER_42_735 VDD VSS sg13g2_decap_8
XFILLER_27_798 VDD VSS sg13g2_decap_8
XFILLER_15_938 VDD VSS sg13g2_decap_8
XFILLER_14_448 VDD VSS sg13g2_decap_8
XFILLER_41_234 VDD VSS sg13g2_decap_8
XFILLER_10_665 VDD VSS sg13g2_decap_8
XFILLER_108_542 VDD VSS sg13g2_decap_8
XFILLER_6_658 VDD VSS sg13g2_decap_8
XFILLER_5_168 VDD VSS sg13g2_decap_8
XFILLER_78_42 VDD VSS sg13g2_decap_8
XFILLER_111_707 VDD VSS sg13g2_decap_8
XFILLER_2_875 VDD VSS sg13g2_decap_8
XFILLER_104_792 VDD VSS sg13g2_decap_8
XFILLER_77_632 VDD VSS sg13g2_decap_8
XFILLER_77_621 VDD VSS sg13g2_decap_4
XFILLER_110_217 VDD VSS sg13g2_decap_8
XFILLER_1_385 VDD VSS sg13g2_decap_8
XFILLER_49_323 VDD VSS sg13g2_decap_8
XFILLER_103_291 VDD VSS sg13g2_decap_8
XFILLER_92_635 VDD VSS sg13g2_fill_2
XFILLER_76_175 VDD VSS sg13g2_decap_8
XFILLER_94_63 VDD VSS sg13g2_decap_8
XFILLER_65_827 VDD VSS sg13g2_decap_8
XFILLER_37_518 VDD VSS sg13g2_decap_8
XFILLER_92_668 VDD VSS sg13g2_decap_8
XFILLER_18_721 VDD VSS sg13g2_decap_8
XFILLER_91_178 VDD VSS sg13g2_decap_4
XFILLER_17_231 VDD VSS sg13g2_decap_8
X_2193__154 VDD VSS _2193_/RESET_B sg13g2_tiehi
XFILLER_33_735 VDD VSS sg13g2_decap_8
XFILLER_60_510 VDD VSS sg13g2_decap_8
XFILLER_18_798 VDD VSS sg13g2_decap_8
XFILLER_32_245 VDD VSS sg13g2_decap_8
XFILLER_60_598 VDD VSS sg13g2_decap_8
XFILLER_41_790 VDD VSS sg13g2_decap_8
XFILLER_9_441 VDD VSS sg13g2_decap_8
X_1514_ _1514_/A _1516_/B _1514_/Y VDD VSS sg13g2_nor2b_1
XFILLER_102_707 VDD VSS sg13g2_decap_8
XFILLER_102_718 VDD VSS sg13g2_fill_2
XFILLER_102_729 VDD VSS sg13g2_fill_2
XFILLER_99_256 VDD VSS sg13g2_decap_8
X_1445_ VDD _2242_/D _1445_/A VSS sg13g2_inv_1
X_1376_ _1376_/Y _1376_/A _1465_/C VDD VSS sg13g2_nand2_1
XFILLER_56_805 VDD VSS sg13g2_decap_8
XFILLER_96_985 VDD VSS sg13g2_decap_8
XFILLER_110_795 VDD VSS sg13g2_decap_8
XFILLER_95_462 VDD VSS sg13g2_decap_8
XFILLER_68_687 VDD VSS sg13g2_decap_8
XFILLER_55_315 VDD VSS sg13g2_decap_8
XFILLER_67_153 VDD VSS sg13g2_decap_8
XFILLER_28_518 VDD VSS sg13g2_decap_8
XFILLER_49_890 VDD VSS sg13g2_decap_8
XFILLER_55_348 VDD VSS sg13g2_decap_8
XFILLER_71_819 VDD VSS sg13g2_decap_8
XFILLER_82_156 VDD VSS sg13g2_decap_8
XFILLER_91_690 VDD VSS sg13g2_decap_8
XFILLER_36_595 VDD VSS sg13g2_decap_8
XFILLER_24_735 VDD VSS sg13g2_decap_8
XFILLER_51_565 VDD VSS sg13g2_decap_8
XFILLER_23_245 VDD VSS sg13g2_decap_8
XFILLER_104_1013 VDD VSS sg13g2_decap_8
XFILLER_17_1043 VDD VSS sg13g2_decap_8
XFILLER_20_952 VDD VSS sg13g2_decap_8
XFILLER_109_306 VDD VSS sg13g2_decap_4
XFILLER_105_512 VDD VSS sg13g2_decap_8
XFILLER_2_105 VDD VSS sg13g2_decap_8
XFILLER_3_7 VDD VSS sg13g2_decap_8
XFILLER_105_567 VDD VSS sg13g2_decap_8
XFILLER_87_941 VDD VSS sg13g2_fill_2
XFILLER_87_963 VDD VSS sg13g2_decap_4
XFILLER_101_740 VDD VSS sg13g2_fill_2
XFILLER_101_751 VDD VSS sg13g2_decap_8
XFILLER_86_440 VDD VSS sg13g2_decap_8
XFILLER_24_1036 VDD VSS sg13g2_decap_8
XFILLER_48_56 VDD VSS sg13g2_decap_8
XFILLER_58_142 VDD VSS sg13g2_decap_8
XFILLER_100_261 VDD VSS sg13g2_decap_8
XFILLER_47_838 VDD VSS sg13g2_decap_8
XFILLER_19_518 VDD VSS sg13g2_decap_8
XFILLER_74_646 VDD VSS sg13g2_decap_8
XFILLER_74_635 VDD VSS sg13g2_fill_1
XFILLER_73_112 VDD VSS sg13g2_decap_8
XFILLER_46_326 VDD VSS sg13g2_decap_8
XFILLER_104_84 VDD VSS sg13g2_decap_8
XFILLER_55_860 VDD VSS sg13g2_decap_8
XFILLER_73_178 VDD VSS sg13g2_decap_8
XFILLER_27_595 VDD VSS sg13g2_decap_8
XFILLER_15_735 VDD VSS sg13g2_decap_8
XFILLER_54_392 VDD VSS sg13g2_fill_1
XFILLER_14_245 VDD VSS sg13g2_decap_8
XFILLER_64_99 VDD VSS sg13g2_decap_8
XFILLER_70_885 VDD VSS sg13g2_decap_8
XFILLER_80_21 VDD VSS sg13g2_decap_8
XFILLER_9_28 VDD VSS sg13g2_decap_8
XFILLER_70_1034 VDD VSS sg13g2_fill_1
Xfanout60 _2270_/Q _2144_/S1 VDD VSS sg13g2_buf_1
XFILLER_30_749 VDD VSS sg13g2_decap_8
XFILLER_11_952 VDD VSS sg13g2_decap_8
Xfanout71 _2107_/B1 _1602_/B VDD VSS sg13g2_buf_1
XFILLER_80_98 VDD VSS sg13g2_decap_8
XFILLER_31_1029 VDD VSS sg13g2_decap_8
XFILLER_10_462 VDD VSS sg13g2_decap_8
XFILLER_109_840 VDD VSS sg13g2_decap_8
XFILLER_13_70 VDD VSS sg13g2_decap_8
XFILLER_7_945 VDD VSS sg13g2_decap_8
X_2223__94 VDD VSS _2223__94/L_HI sg13g2_tiehi
XFILLER_6_455 VDD VSS sg13g2_decap_8
XFILLER_89_63 VDD VSS sg13g2_decap_8
XFILLER_111_504 VDD VSS sg13g2_decap_8
XFILLER_69_407 VDD VSS sg13g2_decap_8
XFILLER_9_1008 VDD VSS sg13g2_decap_8
XFILLER_78_930 VDD VSS sg13g2_decap_8
XFILLER_69_429 VDD VSS sg13g2_fill_2
XFILLER_2_672 VDD VSS sg13g2_decap_8
XFILLER_36_7 VDD VSS sg13g2_decap_8
XFILLER_96_259 VDD VSS sg13g2_decap_8
XFILLER_1_182 VDD VSS sg13g2_decap_8
X_1230_ _1495_/A _1465_/B _1235_/A VDD VSS hold295/X sg13g2_nand3b_1
XFILLER_37_315 VDD VSS sg13g2_decap_8
XFILLER_49_175 VDD VSS sg13g2_decap_8
XFILLER_93_944 VDD VSS sg13g2_decap_8
XFILLER_38_849 VDD VSS sg13g2_decap_8
XFILLER_80_616 VDD VSS sg13g2_decap_8
XFILLER_92_498 VDD VSS sg13g2_decap_8
XFILLER_18_595 VDD VSS sg13g2_decap_8
XFILLER_45_381 VDD VSS sg13g2_decap_8
XFILLER_33_532 VDD VSS sg13g2_decap_8
X_1994_ _1995_/C _1988_/B _1993_/Y _1980_/B _1982_/C VDD VSS sg13g2_a22oi_1
XFILLER_21_749 VDD VSS sg13g2_decap_8
XFILLER_20_259 VDD VSS sg13g2_decap_8
XFILLER_62_0 VDD VSS sg13g2_decap_8
XFILLER_86_1041 VDD VSS sg13g2_decap_8
XFILLER_0_609 VDD VSS sg13g2_decap_8
XFILLER_87_215 VDD VSS sg13g2_fill_2
XFILLER_87_248 VDD VSS sg13g2_decap_8
XFILLER_87_237 VDD VSS sg13g2_fill_2
X_1428_ _2265_/Q _1410_/B _1428_/Y VDD VSS sg13g2_nor2b_1
XFILLER_29_805 VDD VSS sg13g2_decap_8
XFILLER_96_782 VDD VSS sg13g2_decap_8
XFILLER_56_602 VDD VSS sg13g2_decap_8
XFILLER_68_473 VDD VSS sg13g2_decap_8
XFILLER_28_315 VDD VSS sg13g2_decap_8
XFILLER_110_592 VDD VSS sg13g2_decap_8
XFILLER_83_410 VDD VSS sg13g2_decap_8
X_1359_ VDD _2208_/D _1359_/A VSS sg13g2_inv_1
XFILLER_55_123 VDD VSS sg13g2_fill_2
XFILLER_71_605 VDD VSS sg13g2_decap_8
XFILLER_83_487 VDD VSS sg13g2_decap_8
XFILLER_70_126 VDD VSS sg13g2_decap_8
XFILLER_64_690 VDD VSS sg13g2_decap_8
XFILLER_37_882 VDD VSS sg13g2_decap_8
XFILLER_55_189 VDD VSS sg13g2_decap_8
XFILLER_52_863 VDD VSS sg13g2_decap_8
XFILLER_51_340 VDD VSS sg13g2_decap_8
XFILLER_34_14 VDD VSS sg13g2_decap_8
XFILLER_24_532 VDD VSS sg13g2_decap_8
XFILLER_36_392 VDD VSS sg13g2_decap_8
XFILLER_54_1029 VDD VSS sg13g2_decap_8
XFILLER_51_395 VDD VSS sg13g2_decap_8
XFILLER_12_749 VDD VSS sg13g2_decap_8
XFILLER_11_259 VDD VSS sg13g2_decap_8
Xclkload2 VDD clkload2/Y clkload2/A VSS sg13g2_inv_1
XFILLER_109_147 VDD VSS sg13g2_decap_8
XFILLER_50_79 VDD VSS sg13g2_decap_8
XFILLER_106_832 VDD VSS sg13g2_decap_8
XFILLER_4_959 VDD VSS sg13g2_decap_8
XFILLER_3_469 VDD VSS sg13g2_decap_8
XFILLER_105_386 VDD VSS sg13g2_decap_8
XFILLER_75_911 VDD VSS sg13g2_decap_8
XFILLER_93_207 VDD VSS sg13g2_fill_1
XFILLER_75_21 VDD VSS sg13g2_decap_8
XFILLER_47_602 VDD VSS sg13g2_decap_8
XFILLER_86_281 VDD VSS sg13g2_decap_8
XFILLER_86_292 VDD VSS sg13g2_decap_8
XFILLER_74_410 VDD VSS sg13g2_decap_8
XFILLER_19_315 VDD VSS sg13g2_decap_8
XFILLER_75_977 VDD VSS sg13g2_fill_2
XFILLER_75_98 VDD VSS sg13g2_decap_8
XFILLER_35_819 VDD VSS sg13g2_decap_8
XFILLER_46_145 VDD VSS sg13g2_fill_2
XFILLER_62_638 VDD VSS sg13g2_fill_1
XFILLER_28_882 VDD VSS sg13g2_decap_8
XFILLER_61_115 VDD VSS sg13g2_fill_2
XFILLER_34_329 VDD VSS sg13g2_decap_8
XFILLER_46_178 VDD VSS sg13g2_decap_8
XFILLER_91_42 VDD VSS sg13g2_decap_8
XFILLER_43_863 VDD VSS sg13g2_decap_8
XFILLER_15_532 VDD VSS sg13g2_decap_8
XFILLER_27_392 VDD VSS sg13g2_decap_8
XFILLER_70_682 VDD VSS sg13g2_decap_8
XFILLER_30_546 VDD VSS sg13g2_decap_8
XFILLER_42_384 VDD VSS sg13g2_decap_8
XFILLER_24_91 VDD VSS sg13g2_decap_8
XFILLER_7_742 VDD VSS sg13g2_decap_8
XFILLER_6_252 VDD VSS sg13g2_decap_8
X_2331_ _2331_/RESET_B VSS VDD _2331_/D _2331_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_111_301 VDD VSS sg13g2_decap_8
XFILLER_97_513 VDD VSS sg13g2_decap_4
XFILLER_69_204 VDD VSS sg13g2_decap_8
XFILLER_112_868 VDD VSS sg13g2_decap_8
XFILLER_85_708 VDD VSS sg13g2_decap_8
X_2262_ _2262_/RESET_B VSS VDD _2262_/D _2262_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_78_782 VDD VSS sg13g2_decap_8
XFILLER_111_378 VDD VSS sg13g2_decap_8
XFILLER_84_207 VDD VSS sg13g2_decap_8
X_1213_ VDD _1213_/Y _2246_/Q VSS sg13g2_inv_1
XFILLER_66_900 VDD VSS sg13g2_decap_8
X_2193_ _2193_/RESET_B VSS VDD _2193_/D _2193_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_38_646 VDD VSS sg13g2_decap_8
XFILLER_37_112 VDD VSS sg13g2_decap_8
XFILLER_77_1007 VDD VSS sg13g2_decap_8
XFILLER_93_752 VDD VSS sg13g2_decap_8
XFILLER_81_914 VDD VSS sg13g2_decap_4
XFILLER_66_977 VDD VSS sg13g2_decap_8
XFILLER_26_819 VDD VSS sg13g2_decap_8
XFILLER_81_925 VDD VSS sg13g2_decap_8
XFILLER_92_284 VDD VSS sg13g2_fill_2
XFILLER_53_616 VDD VSS sg13g2_decap_8
XFILLER_65_487 VDD VSS sg13g2_decap_8
XFILLER_1_84 VDD VSS sg13g2_decap_8
XFILLER_19_882 VDD VSS sg13g2_decap_8
XFILLER_25_329 VDD VSS sg13g2_decap_8
XFILLER_37_189 VDD VSS sg13g2_decap_8
XFILLER_80_446 VDD VSS sg13g2_decap_8
XFILLER_18_392 VDD VSS sg13g2_decap_8
XFILLER_34_896 VDD VSS sg13g2_decap_8
XFILLER_21_546 VDD VSS sg13g2_decap_8
X_1977_ _2000_/A _1975_/Y _1973_/B _1974_/X _1973_/Y VDD VSS sg13g2_a22oi_1
XFILLER_14_1057 VDD VSS sg13g2_decap_4
XFILLER_101_1016 VDD VSS sg13g2_decap_8
XFILLER_107_618 VDD VSS sg13g2_decap_8
XFILLER_20_49 VDD VSS sg13g2_decap_8
XFILLER_102_312 VDD VSS sg13g2_decap_8
XFILLER_102_301 VDD VSS sg13g2_fill_2
XFILLER_0_406 VDD VSS sg13g2_decap_8
XFILLER_88_568 VDD VSS sg13g2_decap_8
XFILLER_29_14 VDD VSS sg13g2_decap_8
XFILLER_60_1011 VDD VSS sg13g2_decap_8
XFILLER_57_922 VDD VSS sg13g2_decap_8
XFILLER_29_602 VDD VSS sg13g2_decap_8
XFILLER_102_389 VDD VSS sg13g2_decap_8
XFILLER_75_229 VDD VSS sg13g2_decap_8
XFILLER_68_270 VDD VSS sg13g2_decap_8
XFILLER_28_112 VDD VSS sg13g2_decap_8
XFILLER_84_774 VDD VSS sg13g2_decap_8
XFILLER_29_679 VDD VSS sg13g2_decap_8
XFILLER_56_454 VDD VSS sg13g2_decap_8
XFILLER_17_819 VDD VSS sg13g2_decap_8
XFILLER_44_627 VDD VSS sg13g2_decap_8
XFILLER_56_476 VDD VSS sg13g2_decap_8
XFILLER_16_329 VDD VSS sg13g2_decap_8
XFILLER_45_35 VDD VSS sg13g2_decap_8
XFILLER_28_189 VDD VSS sg13g2_decap_8
XFILLER_72_969 VDD VSS sg13g2_decap_8
XFILLER_71_446 VDD VSS sg13g2_decap_8
XFILLER_43_126 VDD VSS sg13g2_decap_8
XFILLER_80_980 VDD VSS sg13g2_decap_8
XFILLER_25_896 VDD VSS sg13g2_decap_8
XFILLER_101_63 VDD VSS sg13g2_decap_8
XFILLER_40_844 VDD VSS sg13g2_decap_8
XFILLER_12_546 VDD VSS sg13g2_decap_8
XFILLER_51_181 VDD VSS sg13g2_decap_8
XFILLER_61_56 VDD VSS sg13g2_decap_8
XFILLER_8_539 VDD VSS sg13g2_decap_8
XFILLER_4_756 VDD VSS sg13g2_decap_8
XFILLER_3_266 VDD VSS sg13g2_decap_8
XFILLER_79_568 VDD VSS sg13g2_decap_4
XFILLER_105_194 VDD VSS sg13g2_decap_8
XFILLER_86_42 VDD VSS sg13g2_decap_8
XFILLER_0_973 VDD VSS sg13g2_decap_8
XFILLER_94_549 VDD VSS sg13g2_decap_8
XFILLER_87_590 VDD VSS sg13g2_decap_8
XFILLER_48_944 VDD VSS sg13g2_decap_8
XFILLER_19_112 VDD VSS sg13g2_decap_8
XFILLER_75_763 VDD VSS sg13g2_fill_1
XFILLER_48_988 VDD VSS sg13g2_decap_8
XFILLER_19_91 VDD VSS sg13g2_decap_8
XFILLER_47_465 VDD VSS sg13g2_fill_2
XFILLER_75_796 VDD VSS sg13g2_decap_4
XFILLER_74_251 VDD VSS sg13g2_decap_8
XFILLER_35_616 VDD VSS sg13g2_decap_8
XFILLER_19_189 VDD VSS sg13g2_decap_8
XFILLER_90_766 VDD VSS sg13g2_decap_8
XFILLER_62_435 VDD VSS sg13g2_decap_8
XFILLER_34_126 VDD VSS sg13g2_decap_8
XFILLER_76_1051 VDD VSS sg13g2_decap_8
XFILLER_90_799 VDD VSS sg13g2_decap_8
XFILLER_43_660 VDD VSS sg13g2_decap_8
XFILLER_71_991 VDD VSS sg13g2_decap_8
X_1900_ _1900_/B _1900_/A _1901_/B VDD VSS sg13g2_xor2_1
XFILLER_37_1057 VDD VSS sg13g2_decap_4
XFILLER_31_833 VDD VSS sg13g2_decap_8
XFILLER_16_896 VDD VSS sg13g2_decap_8
XFILLER_42_170 VDD VSS sg13g2_decap_8
X_1831_ _2249_/Q _2208_/Q _1862_/A VDD VSS sg13g2_nor2b_1
XFILLER_30_343 VDD VSS sg13g2_decap_8
X_1762_ _1762_/B _1762_/A _1888_/A VDD VSS sg13g2_xor2_1
Xhold506 _2316_/Q VDD VSS hold506/X sg13g2_dlygate4sd3_1
Xhold517 _2246_/Q VDD VSS _1453_/A sg13g2_dlygate4sd3_1
X_1693_ _1698_/A _1693_/A _1704_/A VDD VSS sg13g2_xnor2_1
Xhold539 _2318_/Q VDD VSS hold539/X sg13g2_dlygate4sd3_1
Xhold528 _1603_/Y VDD VSS _1604_/B sg13g2_dlygate4sd3_1
XFILLER_97_343 VDD VSS sg13g2_decap_8
XFILLER_112_665 VDD VSS sg13g2_decap_8
XFILLER_98_877 VDD VSS sg13g2_decap_8
X_2314_ _2314_/RESET_B VSS VDD _2314_/D _2314_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_57_207 VDD VSS sg13g2_decap_8
XFILLER_25_0 VDD VSS sg13g2_decap_8
XFILLER_111_175 VDD VSS sg13g2_decap_8
X_2245_ _2245_/RESET_B VSS VDD _2245_/D _2245_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_39_955 VDD VSS sg13g2_decap_8
X_2176_ _2176_/RESET_B VSS VDD _2176_/D _2176_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_65_240 VDD VSS sg13g2_decap_8
XFILLER_38_432 VDD VSS sg13g2_decap_8
XFILLER_93_593 VDD VSS sg13g2_decap_8
XFILLER_81_722 VDD VSS sg13g2_decap_8
XFILLER_26_616 VDD VSS sg13g2_decap_8
XFILLER_65_262 VDD VSS sg13g2_decap_8
XFILLER_54_969 VDD VSS sg13g2_decap_8
XFILLER_20_1050 VDD VSS sg13g2_decap_8
XFILLER_25_126 VDD VSS sg13g2_decap_8
XFILLER_80_276 VDD VSS sg13g2_decap_8
XFILLER_41_608 VDD VSS sg13g2_decap_8
XFILLER_90_1015 VDD VSS sg13g2_decap_8
XFILLER_34_693 VDD VSS sg13g2_decap_8
XFILLER_22_833 VDD VSS sg13g2_decap_8
XFILLER_15_49 VDD VSS sg13g2_decap_8
XFILLER_21_343 VDD VSS sg13g2_decap_8
XFILLER_108_927 VDD VSS sg13g2_decap_8
XFILLER_107_437 VDD VSS sg13g2_decap_8
XFILLER_103_7 VDD VSS sg13g2_decap_8
X_2284__169 VDD VSS _2284_/RESET_B sg13g2_tiehi
XFILLER_0_203 VDD VSS sg13g2_decap_8
XFILLER_89_866 VDD VSS sg13g2_decap_8
XFILLER_88_332 VDD VSS sg13g2_decap_8
XFILLER_103_665 VDD VSS sg13g2_decap_8
XFILLER_76_505 VDD VSS sg13g2_decap_8
XFILLER_102_175 VDD VSS sg13g2_decap_8
XFILLER_88_387 VDD VSS sg13g2_decap_8
XFILLER_57_730 VDD VSS sg13g2_decap_8
XFILLER_5_1022 VDD VSS sg13g2_decap_8
XFILLER_45_947 VDD VSS sg13g2_decap_8
XFILLER_17_616 VDD VSS sg13g2_decap_8
XFILLER_56_67 VDD VSS sg13g2_decap_4
XFILLER_29_476 VDD VSS sg13g2_decap_8
XFILLER_72_766 VDD VSS sg13g2_decap_8
XFILLER_56_284 VDD VSS sg13g2_decap_8
XFILLER_16_126 VDD VSS sg13g2_decap_8
XFILLER_44_446 VDD VSS sg13g2_decap_8
XFILLER_71_276 VDD VSS sg13g2_fill_1
XFILLER_71_265 VDD VSS sg13g2_fill_1
XFILLER_112_84 VDD VSS sg13g2_decap_8
XFILLER_60_928 VDD VSS sg13g2_decap_8
XFILLER_71_287 VDD VSS sg13g2_decap_4
XFILLER_72_77 VDD VSS sg13g2_fill_2
XFILLER_25_693 VDD VSS sg13g2_decap_8
XFILLER_13_833 VDD VSS sg13g2_decap_8
XFILLER_40_641 VDD VSS sg13g2_decap_8
XFILLER_12_343 VDD VSS sg13g2_decap_8
XFILLER_9_826 VDD VSS sg13g2_decap_8
XFILLER_8_336 VDD VSS sg13g2_decap_8
XFILLER_67_1039 VDD VSS sg13g2_decap_8
XFILLER_67_1006 VDD VSS sg13g2_decap_4
XFILLER_21_70 VDD VSS sg13g2_decap_8
XFILLER_107_982 VDD VSS sg13g2_decap_8
XFILLER_106_470 VDD VSS sg13g2_decap_8
XFILLER_4_553 VDD VSS sg13g2_decap_8
XFILLER_97_63 VDD VSS sg13g2_decap_8
XFILLER_95_847 VDD VSS sg13g2_fill_1
XFILLER_95_836 VDD VSS sg13g2_decap_8
XFILLER_79_398 VDD VSS sg13g2_decap_8
XFILLER_0_770 VDD VSS sg13g2_decap_8
X_2030_ _2030_/Y _2074_/A _2030_/B VDD VSS sg13g2_nand2_1
XFILLER_36_903 VDD VSS sg13g2_decap_8
XFILLER_75_560 VDD VSS sg13g2_decap_8
XFILLER_35_413 VDD VSS sg13g2_decap_8
XFILLER_63_744 VDD VSS sg13g2_decap_8
XFILLER_90_563 VDD VSS sg13g2_decap_8
XFILLER_51_939 VDD VSS sg13g2_decap_8
XFILLER_50_416 VDD VSS sg13g2_decap_8
XFILLER_44_991 VDD VSS sg13g2_decap_8
XFILLER_62_287 VDD VSS sg13g2_decap_8
XFILLER_16_693 VDD VSS sg13g2_decap_8
XFILLER_31_630 VDD VSS sg13g2_decap_8
XFILLER_30_140 VDD VSS sg13g2_decap_8
X_1814_ _2219_/Q _2211_/Q _1999_/A VDD VSS sg13g2_xor2_1
XIO_CORNER_NORTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
X_1745_ _2239_/Q _2231_/Q _1763_/B VDD VSS sg13g2_xor2_1
Xhold303 _1276_/Y VDD VSS _1277_/A sg13g2_dlygate4sd3_1
Xhold325 _2165_/Q VDD VSS hold325/X sg13g2_dlygate4sd3_1
Xhold314 _2196_/Q VDD VSS hold314/X sg13g2_dlygate4sd3_1
Xhold358 _1292_/Y VDD VSS _1293_/A sg13g2_dlygate4sd3_1
Xhold369 _1336_/Y VDD VSS _1337_/A sg13g2_dlygate4sd3_1
Xhold336 _2172_/Q VDD VSS hold336/X sg13g2_dlygate4sd3_1
X_1676_ _1680_/B _1677_/A _1677_/B VDD VSS sg13g2_nand2_1
Xhold347 _2357_/Q VDD VSS _2093_/A sg13g2_dlygate4sd3_1
XFILLER_100_602 VDD VSS sg13g2_decap_8
XFILLER_112_462 VDD VSS sg13g2_decap_8
XFILLER_97_151 VDD VSS sg13g2_fill_1
XFILLER_97_140 VDD VSS sg13g2_decap_8
XFILLER_85_313 VDD VSS sg13g2_decap_8
XFILLER_100_668 VDD VSS sg13g2_decap_8
XFILLER_86_869 VDD VSS sg13g2_decap_8
XFILLER_39_752 VDD VSS sg13g2_decap_8
XFILLER_27_903 VDD VSS sg13g2_decap_8
X_2228_ _2228__84/L_HI VSS VDD _2228_/D _2228_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_26_413 VDD VSS sg13g2_decap_8
XFILLER_38_273 VDD VSS sg13g2_decap_8
X_2159_ _2162_/A _2160_/B _2347_/D VDD VSS sg13g2_nor2_1
XFILLER_93_390 VDD VSS sg13g2_decap_8
XFILLER_54_744 VDD VSS sg13g2_decap_8
XFILLER_53_210 VDD VSS sg13g2_fill_1
XFILLER_81_552 VDD VSS sg13g2_decap_8
XFILLER_42_917 VDD VSS sg13g2_decap_8
XFILLER_35_980 VDD VSS sg13g2_decap_8
XFILLER_41_416 VDD VSS sg13g2_decap_8
XFILLER_22_630 VDD VSS sg13g2_decap_8
XFILLER_42_14 VDD VSS sg13g2_decap_8
XFILLER_34_490 VDD VSS sg13g2_decap_8
XFILLER_21_140 VDD VSS sg13g2_decap_8
XFILLER_10_847 VDD VSS sg13g2_decap_8
XFILLER_108_724 VDD VSS sg13g2_decap_8
XFILLER_107_245 VDD VSS sg13g2_decap_8
XFILLER_27_1001 VDD VSS sg13g2_decap_8
XFILLER_104_985 VDD VSS sg13g2_decap_8
XFILLER_89_652 VDD VSS sg13g2_decap_8
XFILLER_103_451 VDD VSS sg13g2_decap_8
XFILLER_107_84 VDD VSS sg13g2_decap_8
XFILLER_88_140 VDD VSS sg13g2_decap_8
XFILLER_1_567 VDD VSS sg13g2_decap_8
XFILLER_89_685 VDD VSS sg13g2_decap_8
XFILLER_76_324 VDD VSS sg13g2_decap_8
XFILLER_76_357 VDD VSS sg13g2_fill_2
XFILLER_18_903 VDD VSS sg13g2_decap_8
XFILLER_67_77 VDD VSS sg13g2_decap_8
XFILLER_85_880 VDD VSS sg13g2_decap_8
XFILLER_85_891 VDD VSS sg13g2_fill_1
XFILLER_91_327 VDD VSS sg13g2_decap_8
XFILLER_17_413 VDD VSS sg13g2_decap_8
XFILLER_29_273 VDD VSS sg13g2_decap_8
XFILLER_83_21 VDD VSS sg13g2_decap_8
XFILLER_45_744 VDD VSS sg13g2_decap_8
XFILLER_44_232 VDD VSS sg13g2_fill_2
XFILLER_33_917 VDD VSS sg13g2_decap_8
XFILLER_44_265 VDD VSS sg13g2_decap_8
XFILLER_83_98 VDD VSS sg13g2_decap_8
XFILLER_26_980 VDD VSS sg13g2_decap_8
XFILLER_60_736 VDD VSS sg13g2_decap_8
XFILLER_16_70 VDD VSS sg13g2_decap_8
XFILLER_32_427 VDD VSS sg13g2_decap_8
XFILLER_44_287 VDD VSS sg13g2_decap_8
XFILLER_13_630 VDD VSS sg13g2_decap_8
XFILLER_25_490 VDD VSS sg13g2_decap_8
XFILLER_41_972 VDD VSS sg13g2_decap_8
XFILLER_12_140 VDD VSS sg13g2_decap_8
XFILLER_9_623 VDD VSS sg13g2_decap_8
XFILLER_8_133 VDD VSS sg13g2_decap_8
XFILLER_32_91 VDD VSS sg13g2_decap_8
XFILLER_66_7 VDD VSS sg13g2_decap_8
XFILLER_5_840 VDD VSS sg13g2_decap_8
X_1530_ VSS VDD _1556_/S0 _1215_/Y _1530_/Y _1523_/B sg13g2_a21oi_1
XFILLER_4_350 VDD VSS sg13g2_decap_8
X_1461_ _1461_/A _1463_/B _1461_/Y VDD VSS sg13g2_nor2_1
XFILLER_110_900 VDD VSS sg13g2_decap_8
X_1392_ _1429_/A _1392_/B _1392_/Y VDD VSS sg13g2_nor2_1
XFILLER_79_140 VDD VSS sg13g2_decap_8
XFILLER_110_977 VDD VSS sg13g2_decap_8
XFILLER_68_869 VDD VSS sg13g2_decap_8
XFILLER_67_357 VDD VSS sg13g2_decap_8
XFILLER_55_508 VDD VSS sg13g2_decap_8
XFILLER_94_154 VDD VSS sg13g2_decap_8
XFILLER_36_700 VDD VSS sg13g2_decap_8
X_2013_ _1999_/A _1931_/A _2021_/S _2015_/B VDD VSS sg13g2_mux2_1
XFILLER_82_349 VDD VSS sg13g2_decap_8
XFILLER_48_582 VDD VSS sg13g2_decap_8
XFILLER_35_210 VDD VSS sg13g2_decap_8
XFILLER_24_917 VDD VSS sg13g2_decap_8
XFILLER_63_552 VDD VSS sg13g2_decap_8
XFILLER_51_703 VDD VSS sg13g2_decap_8
XFILLER_36_777 VDD VSS sg13g2_decap_8
XFILLER_90_393 VDD VSS sg13g2_decap_4
XFILLER_17_980 VDD VSS sg13g2_decap_8
XFILLER_23_427 VDD VSS sg13g2_decap_8
XFILLER_35_287 VDD VSS sg13g2_decap_8
XFILLER_50_202 VDD VSS sg13g2_decap_8
XFILLER_92_0 VDD VSS sg13g2_decap_8
XFILLER_51_758 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_15_clk clkbuf_2_2__f_clk/X _2365_/CLK VDD VSS sg13g2_buf_8
XFILLER_16_490 VDD VSS sg13g2_decap_8
XFILLER_32_994 VDD VSS sg13g2_decap_8
XFILLER_12_28 VDD VSS sg13g2_decap_8
XFILLER_89_1050 VDD VSS sg13g2_decap_8
X_1728_ _2230_/Q _2238_/Q _1728_/Y VDD VSS sg13g2_nor2b_1
XFILLER_105_749 VDD VSS sg13g2_decap_8
X_1659_ _2310_/Q _2332_/Q _2324_/Q _2347_/Q _2339_/Q _2311_/Q _1659_/X VDD VSS sg13g2_mux4_1
XFILLER_99_972 VDD VSS sg13g2_decap_8
XFILLER_101_900 VDD VSS sg13g2_decap_8
XFILLER_104_259 VDD VSS sg13g2_decap_8
XFILLER_59_803 VDD VSS sg13g2_decap_8
XFILLER_86_611 VDD VSS sg13g2_fill_2
XFILLER_58_302 VDD VSS sg13g2_decap_8
XFILLER_101_977 VDD VSS sg13g2_decap_8
XFILLER_100_443 VDD VSS sg13g2_fill_1
XFILLER_100_432 VDD VSS sg13g2_decap_8
XFILLER_85_143 VDD VSS sg13g2_decap_8
XFILLER_37_14 VDD VSS sg13g2_decap_8
XFILLER_74_828 VDD VSS sg13g2_decap_8
XFILLER_27_700 VDD VSS sg13g2_decap_8
XFILLER_96_1032 VDD VSS sg13g2_decap_8
XFILLER_2_1036 VDD VSS sg13g2_decap_8
XFILLER_26_210 VDD VSS sg13g2_decap_8
XFILLER_82_872 VDD VSS sg13g2_decap_8
XFILLER_42_714 VDD VSS sg13g2_decap_8
XFILLER_27_777 VDD VSS sg13g2_decap_8
XFILLER_15_917 VDD VSS sg13g2_decap_8
XFILLER_14_427 VDD VSS sg13g2_decap_8
XFILLER_26_287 VDD VSS sg13g2_decap_8
XFILLER_41_202 VDD VSS sg13g2_decap_8
XFILLER_23_994 VDD VSS sg13g2_decap_8
XFILLER_50_791 VDD VSS sg13g2_decap_8
XFILLER_10_644 VDD VSS sg13g2_decap_8
XFILLER_108_521 VDD VSS sg13g2_decap_8
XFILLER_6_637 VDD VSS sg13g2_decap_8
XFILLER_5_147 VDD VSS sg13g2_decap_8
XFILLER_108_598 VDD VSS sg13g2_decap_8
XFILLER_97_909 VDD VSS sg13g2_decap_8
XFILLER_78_21 VDD VSS sg13g2_decap_8
XFILLER_64_1009 VDD VSS sg13g2_fill_1
XFILLER_2_854 VDD VSS sg13g2_decap_8
XFILLER_104_771 VDD VSS sg13g2_decap_8
XFILLER_77_600 VDD VSS sg13g2_decap_8
XFILLER_103_270 VDD VSS sg13g2_decap_8
XFILLER_78_98 VDD VSS sg13g2_decap_8
XFILLER_1_364 VDD VSS sg13g2_decap_8
XFILLER_49_302 VDD VSS sg13g2_decap_8
XFILLER_65_806 VDD VSS sg13g2_decap_8
XFILLER_92_614 VDD VSS sg13g2_decap_8
XFILLER_77_688 VDD VSS sg13g2_decap_8
XFILLER_94_42 VDD VSS sg13g2_decap_8
XFILLER_76_154 VDD VSS sg13g2_decap_8
XFILLER_18_700 VDD VSS sg13g2_decap_8
XFILLER_92_647 VDD VSS sg13g2_decap_8
XFILLER_57_390 VDD VSS sg13g2_decap_8
XFILLER_17_210 VDD VSS sg13g2_decap_8
XFILLER_91_157 VDD VSS sg13g2_decap_8
XFILLER_18_777 VDD VSS sg13g2_decap_8
XFILLER_73_894 VDD VSS sg13g2_decap_8
XFILLER_45_574 VDD VSS sg13g2_decap_8
XFILLER_33_714 VDD VSS sg13g2_decap_8
XFILLER_17_287 VDD VSS sg13g2_decap_8
XFILLER_27_91 VDD VSS sg13g2_decap_8
XFILLER_60_566 VDD VSS sg13g2_decap_8
XFILLER_32_224 VDD VSS sg13g2_decap_8
XFILLER_14_994 VDD VSS sg13g2_decap_8
X_2269__215 VDD VSS _2269_/RESET_B sg13g2_tiehi
XFILLER_9_420 VDD VSS sg13g2_decap_8
XFILLER_9_497 VDD VSS sg13g2_decap_8
XFILLER_99_235 VDD VSS sg13g2_decap_8
XFILLER_99_213 VDD VSS sg13g2_fill_2
X_1513_ _1671_/C _1513_/B _1513_/C _1513_/Y VDD VSS sg13g2_nor3_1
XFILLER_96_920 VDD VSS sg13g2_decap_8
X_1444_ _1445_/A _1429_/Y hold536/X _1428_/Y _1388_/A VDD VSS sg13g2_a22oi_1
Xclkbuf_leaf_4_clk clkbuf_leaf_5_clk/A clkload6/A VDD VSS sg13g2_buf_8
XFILLER_68_622 VDD VSS sg13g2_decap_8
XFILLER_4_84 VDD VSS sg13g2_decap_8
X_2280__183 VDD VSS _2280_/RESET_B sg13g2_tiehi
XFILLER_95_441 VDD VSS sg13g2_decap_8
X_1375_ _1374_/Y VDD _2213_/D VSS _1367_/B _1373_/Y sg13g2_o21ai_1
XFILLER_68_666 VDD VSS sg13g2_decap_8
XFILLER_110_774 VDD VSS sg13g2_decap_8
XFILLER_83_647 VDD VSS sg13g2_decap_8
XFILLER_64_894 VDD VSS sg13g2_decap_8
XFILLER_36_574 VDD VSS sg13g2_decap_8
XFILLER_24_714 VDD VSS sg13g2_decap_8
XFILLER_51_544 VDD VSS sg13g2_decap_8
XFILLER_23_224 VDD VSS sg13g2_decap_8
XFILLER_17_1022 VDD VSS sg13g2_decap_8
XFILLER_32_791 VDD VSS sg13g2_decap_8
XFILLER_20_931 VDD VSS sg13g2_decap_8
XFILLER_23_49 VDD VSS sg13g2_decap_8
XFILLER_99_780 VDD VSS sg13g2_decap_8
XFILLER_24_1015 VDD VSS sg13g2_decap_8
XFILLER_59_644 VDD VSS sg13g2_decap_8
XFILLER_48_35 VDD VSS sg13g2_decap_8
XFILLER_58_121 VDD VSS sg13g2_decap_8
XFILLER_87_997 VDD VSS sg13g2_decap_8
XFILLER_100_240 VDD VSS sg13g2_decap_8
XFILLER_47_817 VDD VSS sg13g2_decap_8
XFILLER_111_1029 VDD VSS sg13g2_decap_8
XFILLER_86_496 VDD VSS sg13g2_fill_1
XFILLER_104_63 VDD VSS sg13g2_decap_8
XFILLER_58_187 VDD VSS sg13g2_decap_8
XFILLER_73_157 VDD VSS sg13g2_decap_8
XFILLER_27_574 VDD VSS sg13g2_decap_8
XFILLER_15_714 VDD VSS sg13g2_decap_8
XFILLER_64_56 VDD VSS sg13g2_decap_8
XFILLER_70_864 VDD VSS sg13g2_decap_8
XFILLER_14_224 VDD VSS sg13g2_decap_8
XFILLER_42_588 VDD VSS sg13g2_decap_8
XFILLER_30_728 VDD VSS sg13g2_decap_8
Xfanout72 _2107_/B1 _1367_/A VDD VSS sg13g2_buf_1
Xfanout61 _2124_/A _1510_/A VDD VSS sg13g2_buf_1
XFILLER_23_791 VDD VSS sg13g2_decap_8
XFILLER_11_931 VDD VSS sg13g2_decap_8
Xfanout50 _2288_/Q _1592_/A VDD VSS sg13g2_buf_1
XFILLER_80_77 VDD VSS sg13g2_decap_8
XFILLER_31_1008 VDD VSS sg13g2_decap_8
XFILLER_10_441 VDD VSS sg13g2_decap_8
XFILLER_7_924 VDD VSS sg13g2_decap_8
XFILLER_6_434 VDD VSS sg13g2_decap_8
XFILLER_108_340 VDD VSS sg13g2_decap_8
XFILLER_89_42 VDD VSS sg13g2_decap_8
XFILLER_109_896 VDD VSS sg13g2_decap_8
XFILLER_2_651 VDD VSS sg13g2_decap_8
XFILLER_1_161 VDD VSS sg13g2_decap_8
XFILLER_96_238 VDD VSS sg13g2_decap_8
XFILLER_77_430 VDD VSS sg13g2_fill_1
XFILLER_29_7 VDD VSS sg13g2_decap_8
XFILLER_78_986 VDD VSS sg13g2_decap_8
XFILLER_93_901 VDD VSS sg13g2_decap_8
XFILLER_38_828 VDD VSS sg13g2_decap_8
XFILLER_49_154 VDD VSS sg13g2_decap_8
XFILLER_92_422 VDD VSS sg13g2_decap_4
XFILLER_65_658 VDD VSS sg13g2_decap_8
XFILLER_64_113 VDD VSS sg13g2_decap_4
XFILLER_92_477 VDD VSS sg13g2_decap_8
XFILLER_92_455 VDD VSS sg13g2_decap_8
XFILLER_65_669 VDD VSS sg13g2_fill_2
XFILLER_64_157 VDD VSS sg13g2_decap_8
XFILLER_46_894 VDD VSS sg13g2_fill_1
XFILLER_18_574 VDD VSS sg13g2_decap_8
XFILLER_33_511 VDD VSS sg13g2_decap_8
XFILLER_61_886 VDD VSS sg13g2_decap_8
XFILLER_33_588 VDD VSS sg13g2_decap_8
XFILLER_21_728 VDD VSS sg13g2_decap_8
XFILLER_60_352 VDD VSS sg13g2_decap_8
X_1993_ _1993_/Y _2005_/C _1984_/B VDD VSS sg13g2_nand2b_1
XFILLER_20_238 VDD VSS sg13g2_decap_8
XFILLER_14_791 VDD VSS sg13g2_decap_8
XFILLER_9_294 VDD VSS sg13g2_decap_8
XFILLER_55_0 VDD VSS sg13g2_decap_8
X_2323__220 VDD VSS _2323_/RESET_B sg13g2_tiehi
XFILLER_102_505 VDD VSS sg13g2_decap_4
XFILLER_47_1059 VDD VSS sg13g2_fill_2
XFILLER_47_1048 VDD VSS sg13g2_decap_8
X_2362__280 VDD VSS _2362_/RESET_B sg13g2_tiehi
XFILLER_69_964 VDD VSS sg13g2_decap_8
XFILLER_102_549 VDD VSS sg13g2_decap_4
X_1427_ _1426_/Y VDD _2234_/D VSS _1388_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_68_441 VDD VSS sg13g2_fill_2
XFILLER_69_997 VDD VSS sg13g2_fill_1
XFILLER_96_761 VDD VSS sg13g2_decap_8
XFILLER_110_571 VDD VSS sg13g2_decap_8
XFILLER_95_293 VDD VSS sg13g2_decap_8
X_1358_ _1359_/A _1347_/Y hold421/X _1347_/B _1382_/A VDD VSS sg13g2_a22oi_1
XFILLER_18_49 VDD VSS sg13g2_decap_8
XFILLER_55_102 VDD VSS sg13g2_decap_8
XFILLER_110_1040 VDD VSS sg13g2_decap_8
X_1289_ VDD _2174_/D _1289_/A VSS sg13g2_inv_1
XFILLER_83_466 VDD VSS sg13g2_decap_8
XFILLER_56_658 VDD VSS sg13g2_decap_8
XFILLER_37_861 VDD VSS sg13g2_decap_8
XFILLER_43_308 VDD VSS sg13g2_fill_1
XFILLER_70_105 VDD VSS sg13g2_decap_8
XFILLER_55_168 VDD VSS sg13g2_decap_8
XFILLER_24_511 VDD VSS sg13g2_decap_8
XFILLER_36_371 VDD VSS sg13g2_decap_8
XFILLER_52_831 VDD VSS sg13g2_decap_8
XFILLER_54_1019 VDD VSS sg13g2_decap_4
XFILLER_24_588 VDD VSS sg13g2_decap_8
XFILLER_12_728 VDD VSS sg13g2_decap_8
XFILLER_11_238 VDD VSS sg13g2_decap_8
Xclkload3 clkload3/A clkload3/Y VDD VSS sg13g2_inv_4
XFILLER_50_14 VDD VSS sg13g2_decap_8
XFILLER_109_126 VDD VSS sg13g2_decap_8
XFILLER_50_58 VDD VSS sg13g2_decap_8
XFILLER_106_811 VDD VSS sg13g2_decap_8
XFILLER_4_938 VDD VSS sg13g2_decap_8
X_2328__197 VDD VSS _2328_/RESET_B sg13g2_tiehi
XFILLER_3_448 VDD VSS sg13g2_decap_8
XFILLER_106_888 VDD VSS sg13g2_decap_8
XFILLER_105_365 VDD VSS sg13g2_decap_8
XFILLER_75_956 VDD VSS sg13g2_decap_8
XFILLER_87_794 VDD VSS sg13g2_decap_8
XFILLER_46_102 VDD VSS sg13g2_fill_1
XFILLER_46_124 VDD VSS sg13g2_decap_8
XFILLER_75_77 VDD VSS sg13g2_decap_8
XFILLER_47_658 VDD VSS sg13g2_decap_4
XFILLER_28_861 VDD VSS sg13g2_decap_8
XFILLER_90_937 VDD VSS sg13g2_decap_8
XFILLER_62_617 VDD VSS sg13g2_decap_8
XFILLER_15_511 VDD VSS sg13g2_decap_8
XFILLER_27_371 VDD VSS sg13g2_decap_8
XFILLER_34_308 VDD VSS sg13g2_decap_8
XFILLER_91_21 VDD VSS sg13g2_decap_8
XFILLER_43_842 VDD VSS sg13g2_decap_8
XFILLER_70_661 VDD VSS sg13g2_decap_8
XFILLER_15_588 VDD VSS sg13g2_decap_8
XFILLER_42_363 VDD VSS sg13g2_decap_8
XFILLER_91_98 VDD VSS sg13g2_decap_8
XFILLER_30_525 VDD VSS sg13g2_decap_8
XFILLER_24_70 VDD VSS sg13g2_decap_8
XFILLER_7_721 VDD VSS sg13g2_decap_8
XFILLER_6_231 VDD VSS sg13g2_decap_8
XFILLER_109_693 VDD VSS sg13g2_decap_8
XFILLER_7_798 VDD VSS sg13g2_decap_8
XFILLER_40_91 VDD VSS sg13g2_decap_8
X_2330_ _2330_/RESET_B VSS VDD _2330_/D _2330_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_112_847 VDD VSS sg13g2_decap_8
X_2261_ _2261_/RESET_B VSS VDD _2261_/D _2261_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_78_761 VDD VSS sg13g2_decap_8
XFILLER_111_357 VDD VSS sg13g2_decap_8
X_1212_ VDD _1212_/Y _2247_/Q VSS sg13g2_inv_1
X_2192_ _2192_/RESET_B VSS VDD _2192_/D _2192_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_93_731 VDD VSS sg13g2_decap_8
XFILLER_77_260 VDD VSS sg13g2_fill_1
XFILLER_66_956 VDD VSS sg13g2_decap_8
XFILLER_38_625 VDD VSS sg13g2_decap_8
XFILLER_65_466 VDD VSS sg13g2_decap_8
XFILLER_1_63 VDD VSS sg13g2_decap_8
XFILLER_19_861 VDD VSS sg13g2_decap_8
XFILLER_92_263 VDD VSS sg13g2_decap_8
XFILLER_80_425 VDD VSS sg13g2_decap_8
XFILLER_18_371 VDD VSS sg13g2_decap_8
XFILLER_25_308 VDD VSS sg13g2_decap_8
XFILLER_37_168 VDD VSS sg13g2_decap_8
XFILLER_52_138 VDD VSS sg13g2_decap_8
XFILLER_34_875 VDD VSS sg13g2_decap_8
XFILLER_21_525 VDD VSS sg13g2_decap_8
XFILLER_33_385 VDD VSS sg13g2_decap_8
X_1976_ _1976_/Y _1976_/A _1976_/B VDD VSS sg13g2_xnor2_1
XFILLER_60_193 VDD VSS sg13g2_decap_8
XFILLER_14_1036 VDD VSS sg13g2_decap_8
XFILLER_101_1006 VDD VSS sg13g2_fill_1
XFILLER_20_28 VDD VSS sg13g2_decap_8
X_2208__124 VDD VSS _2208_/RESET_B sg13g2_tiehi
XFILLER_103_836 VDD VSS sg13g2_fill_2
XFILLER_88_503 VDD VSS sg13g2_decap_8
XFILLER_88_547 VDD VSS sg13g2_decap_8
XFILLER_102_368 VDD VSS sg13g2_decap_8
XFILLER_75_208 VDD VSS sg13g2_decap_8
XFILLER_57_901 VDD VSS sg13g2_decap_8
XFILLER_69_783 VDD VSS sg13g2_decap_8
XFILLER_68_260 VDD VSS sg13g2_decap_4
XFILLER_57_967 VDD VSS sg13g2_fill_2
XFILLER_21_1029 VDD VSS sg13g2_decap_8
XFILLER_44_606 VDD VSS sg13g2_decap_8
XFILLER_29_658 VDD VSS sg13g2_decap_8
XFILLER_56_433 VDD VSS sg13g2_decap_8
XFILLER_72_948 VDD VSS sg13g2_decap_8
XFILLER_72_937 VDD VSS sg13g2_fill_2
XFILLER_84_797 VDD VSS sg13g2_decap_4
XFILLER_83_285 VDD VSS sg13g2_decap_8
XFILLER_71_425 VDD VSS sg13g2_decap_8
XFILLER_16_308 VDD VSS sg13g2_decap_8
XFILLER_43_105 VDD VSS sg13g2_decap_8
XFILLER_45_14 VDD VSS sg13g2_decap_8
XFILLER_28_168 VDD VSS sg13g2_decap_8
XFILLER_101_42 VDD VSS sg13g2_decap_8
XFILLER_52_661 VDD VSS sg13g2_decap_4
XFILLER_25_875 VDD VSS sg13g2_decap_8
XFILLER_40_823 VDD VSS sg13g2_decap_8
XFILLER_12_525 VDD VSS sg13g2_decap_8
XFILLER_24_385 VDD VSS sg13g2_decap_8
XFILLER_8_518 VDD VSS sg13g2_decap_8
XFILLER_61_35 VDD VSS sg13g2_decap_8
XFILLER_4_735 VDD VSS sg13g2_decap_8
XFILLER_3_245 VDD VSS sg13g2_decap_8
XFILLER_106_685 VDD VSS sg13g2_decap_8
XFILLER_105_140 VDD VSS sg13g2_decap_8
XFILLER_79_547 VDD VSS sg13g2_decap_8
XFILLER_86_21 VDD VSS sg13g2_decap_8
XFILLER_48_901 VDD VSS sg13g2_decap_8
XFILLER_0_952 VDD VSS sg13g2_decap_8
XFILLER_48_923 VDD VSS sg13g2_decap_8
XFILLER_75_742 VDD VSS sg13g2_decap_8
XFILLER_74_230 VDD VSS sg13g2_decap_8
XFILLER_48_956 VDD VSS sg13g2_decap_4
XFILLER_48_967 VDD VSS sg13g2_decap_8
XFILLER_19_70 VDD VSS sg13g2_decap_8
XFILLER_47_455 VDD VSS sg13g2_fill_1
XFILLER_75_775 VDD VSS sg13g2_decap_8
XFILLER_62_414 VDD VSS sg13g2_decap_8
XFILLER_19_168 VDD VSS sg13g2_decap_8
XFILLER_34_105 VDD VSS sg13g2_decap_8
XFILLER_47_488 VDD VSS sg13g2_decap_8
XFILLER_90_745 VDD VSS sg13g2_decap_8
X_2272__211 VDD VSS _2272_/RESET_B sg13g2_tiehi
XFILLER_71_970 VDD VSS sg13g2_decap_8
XFILLER_31_812 VDD VSS sg13g2_decap_8
XFILLER_16_875 VDD VSS sg13g2_decap_8
XFILLER_70_491 VDD VSS sg13g2_decap_8
XFILLER_96_7 VDD VSS sg13g2_decap_8
XFILLER_37_1036 VDD VSS sg13g2_decap_8
XFILLER_15_385 VDD VSS sg13g2_decap_8
XFILLER_35_91 VDD VSS sg13g2_decap_8
XFILLER_30_322 VDD VSS sg13g2_decap_8
X_1830_ _1852_/A _2250_/Q _2209_/Q VDD VSS sg13g2_xnor2_1
XFILLER_31_889 VDD VSS sg13g2_decap_8
X_1761_ _1762_/B _1761_/A _1761_/B VDD VSS sg13g2_nand2_1
XFILLER_30_399 VDD VSS sg13g2_decap_8
Xhold507 _1707_/Y VDD VSS _2316_/D sg13g2_dlygate4sd3_1
X_1692_ _1704_/A _1692_/A _1692_/B VDD VSS sg13g2_xnor2_1
Xhold518 _2262_/Q VDD VSS hold518/X sg13g2_dlygate4sd3_1
XFILLER_109_490 VDD VSS sg13g2_decap_8
XFILLER_7_595 VDD VSS sg13g2_decap_8
Xhold529 _1604_/Y VDD VSS _2290_/D sg13g2_dlygate4sd3_1
XFILLER_83_1012 VDD VSS sg13g2_fill_1
XFILLER_98_834 VDD VSS sg13g2_decap_8
XFILLER_83_1045 VDD VSS sg13g2_decap_8
XFILLER_112_644 VDD VSS sg13g2_decap_8
XFILLER_97_322 VDD VSS sg13g2_decap_8
X_2313_ _2313_/RESET_B VSS VDD _2313_/D _2313_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_111_154 VDD VSS sg13g2_decap_8
X_2244_ _2244_/RESET_B VSS VDD _2244_/D _2244_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_934 VDD VSS sg13g2_decap_8
XFILLER_38_411 VDD VSS sg13g2_decap_8
X_2175_ _2175_/RESET_B VSS VDD _2175_/D _2175_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_18_0 VDD VSS sg13g2_decap_8
XFILLER_93_572 VDD VSS sg13g2_decap_8
XFILLER_81_701 VDD VSS sg13g2_decap_8
XFILLER_54_948 VDD VSS sg13g2_decap_8
XFILLER_66_775 VDD VSS sg13g2_fill_2
XFILLER_53_414 VDD VSS sg13g2_fill_1
XFILLER_53_403 VDD VSS sg13g2_fill_2
XFILLER_25_105 VDD VSS sg13g2_decap_8
XFILLER_38_488 VDD VSS sg13g2_decap_8
XFILLER_81_789 VDD VSS sg13g2_decap_4
XFILLER_80_255 VDD VSS sg13g2_decap_8
XFILLER_15_28 VDD VSS sg13g2_decap_8
XFILLER_62_992 VDD VSS sg13g2_decap_8
XFILLER_34_672 VDD VSS sg13g2_decap_8
XFILLER_22_812 VDD VSS sg13g2_decap_8
XFILLER_40_119 VDD VSS sg13g2_decap_8
XFILLER_21_322 VDD VSS sg13g2_decap_8
XFILLER_33_182 VDD VSS sg13g2_decap_8
XFILLER_22_889 VDD VSS sg13g2_decap_8
XFILLER_108_906 VDD VSS sg13g2_decap_8
X_1959_ _1950_/Y VDD _1962_/A VSS _1955_/A _1955_/B sg13g2_o21ai_1
XFILLER_31_49 VDD VSS sg13g2_decap_8
XFILLER_21_399 VDD VSS sg13g2_decap_8
XFILLER_107_416 VDD VSS sg13g2_decap_8
XFILLER_103_644 VDD VSS sg13g2_decap_8
XFILLER_1_749 VDD VSS sg13g2_decap_8
XFILLER_102_154 VDD VSS sg13g2_decap_8
XFILLER_0_259 VDD VSS sg13g2_decap_8
XFILLER_5_1001 VDD VSS sg13g2_decap_8
XFILLER_102_198 VDD VSS sg13g2_decap_8
XFILLER_29_455 VDD VSS sg13g2_decap_8
XFILLER_45_926 VDD VSS sg13g2_decap_8
XFILLER_57_786 VDD VSS sg13g2_decap_8
XFILLER_56_263 VDD VSS sg13g2_decap_8
XFILLER_16_105 VDD VSS sg13g2_decap_8
XFILLER_44_403 VDD VSS sg13g2_fill_2
XFILLER_72_756 VDD VSS sg13g2_fill_1
X_2256__239 VDD VSS _2256_/RESET_B sg13g2_tiehi
XFILLER_112_63 VDD VSS sg13g2_decap_8
XFILLER_60_907 VDD VSS sg13g2_decap_8
XFILLER_32_609 VDD VSS sg13g2_decap_8
XFILLER_71_299 VDD VSS sg13g2_decap_4
XFILLER_72_56 VDD VSS sg13g2_decap_8
XFILLER_40_620 VDD VSS sg13g2_decap_8
XFILLER_25_672 VDD VSS sg13g2_decap_8
XFILLER_13_812 VDD VSS sg13g2_decap_8
XFILLER_31_119 VDD VSS sg13g2_decap_8
XFILLER_12_322 VDD VSS sg13g2_decap_8
XFILLER_9_805 VDD VSS sg13g2_decap_8
XFILLER_24_182 VDD VSS sg13g2_decap_8
XFILLER_40_697 VDD VSS sg13g2_decap_8
XFILLER_8_315 VDD VSS sg13g2_decap_8
XFILLER_13_889 VDD VSS sg13g2_decap_8
XFILLER_12_399 VDD VSS sg13g2_decap_8
XFILLER_4_532 VDD VSS sg13g2_decap_8
XFILLER_107_961 VDD VSS sg13g2_decap_8
XFILLER_98_119 VDD VSS sg13g2_decap_8
XFILLER_97_42 VDD VSS sg13g2_decap_8
XFILLER_95_815 VDD VSS sg13g2_decap_8
XFILLER_79_355 VDD VSS sg13g2_decap_4
XFILLER_94_303 VDD VSS sg13g2_decap_8
XFILLER_79_377 VDD VSS sg13g2_decap_8
XFILLER_67_539 VDD VSS sg13g2_decap_8
XFILLER_11_7 VDD VSS sg13g2_decap_8
XFILLER_63_723 VDD VSS sg13g2_decap_8
XFILLER_48_775 VDD VSS sg13g2_decap_8
XFILLER_90_542 VDD VSS sg13g2_decap_8
XFILLER_36_959 VDD VSS sg13g2_decap_8
XFILLER_47_285 VDD VSS sg13g2_decap_8
XFILLER_51_918 VDD VSS sg13g2_decap_8
XFILLER_44_970 VDD VSS sg13g2_decap_8
XFILLER_23_609 VDD VSS sg13g2_decap_8
XFILLER_35_469 VDD VSS sg13g2_decap_8
XFILLER_16_672 VDD VSS sg13g2_decap_8
XFILLER_22_119 VDD VSS sg13g2_decap_8
Xclkbuf_0_clk clkbuf_0_clk/X clk_pad/p2c VDD VSS sg13g2_buf_16
XFILLER_15_182 VDD VSS sg13g2_decap_8
XFILLER_31_686 VDD VSS sg13g2_decap_8
X_1813_ _1939_/B _2211_/Q _2219_/Q VDD VSS sg13g2_xnor2_1
XFILLER_30_196 VDD VSS sg13g2_decap_8
X_1744_ _1761_/A _2239_/Q _2231_/Q VDD VSS sg13g2_nand2b_1
XFILLER_8_882 VDD VSS sg13g2_decap_8
Xhold326 _1270_/Y VDD VSS _1271_/A sg13g2_dlygate4sd3_1
Xhold304 _2191_/Q VDD VSS hold304/X sg13g2_dlygate4sd3_1
Xhold315 _1332_/Y VDD VSS _1333_/A sg13g2_dlygate4sd3_1
XFILLER_7_392 VDD VSS sg13g2_decap_8
XFILLER_7_84 VDD VSS sg13g2_decap_8
XFILLER_104_419 VDD VSS sg13g2_fill_2
XFILLER_89_119 VDD VSS sg13g2_decap_8
Xhold337 _1284_/Y VDD VSS _1285_/A sg13g2_dlygate4sd3_1
X_1675_ _1681_/A _1675_/B _1677_/B _1675_/Y VDD VSS sg13g2_nor3_1
Xhold348 _1222_/Y VDD VSS _2363_/D sg13g2_dlygate4sd3_1
Xhold359 _2257_/Q VDD VSS _1196_/A sg13g2_dlygate4sd3_1
XFILLER_98_642 VDD VSS sg13g2_fill_1
XFILLER_112_441 VDD VSS sg13g2_decap_8
XFILLER_98_697 VDD VSS sg13g2_decap_8
XFILLER_86_848 VDD VSS sg13g2_decap_8
XFILLER_86_837 VDD VSS sg13g2_decap_8
X_2227_ _2227__86/L_HI VSS VDD _2227_/D _2227_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_39_731 VDD VSS sg13g2_decap_8
XFILLER_85_369 VDD VSS sg13g2_decap_8
XFILLER_66_561 VDD VSS sg13g2_decap_8
XFILLER_54_712 VDD VSS sg13g2_decap_8
XFILLER_38_252 VDD VSS sg13g2_decap_8
XFILLER_94_892 VDD VSS sg13g2_decap_8
X_2158_ _2162_/A _2162_/B _2346_/D VDD VSS sg13g2_nor2_1
XFILLER_81_531 VDD VSS sg13g2_decap_8
XFILLER_27_959 VDD VSS sg13g2_decap_8
XFILLER_54_723 VDD VSS sg13g2_fill_2
X_2089_ _2068_/B _2071_/C _2089_/S _2149_/B VDD VSS sg13g2_mux2_1
XFILLER_14_609 VDD VSS sg13g2_decap_8
XFILLER_26_49 VDD VSS sg13g2_decap_8
XFILLER_26_469 VDD VSS sg13g2_decap_8
XFILLER_53_299 VDD VSS sg13g2_decap_8
XFILLER_13_119 VDD VSS sg13g2_decap_8
XFILLER_107_1045 VDD VSS sg13g2_decap_8
XFILLER_50_995 VDD VSS sg13g2_decap_8
XFILLER_22_686 VDD VSS sg13g2_decap_8
XFILLER_10_826 VDD VSS sg13g2_decap_8
XFILLER_6_819 VDD VSS sg13g2_decap_8
XFILLER_21_196 VDD VSS sg13g2_decap_8
XFILLER_108_703 VDD VSS sg13g2_decap_8
XFILLER_5_329 VDD VSS sg13g2_decap_8
XFILLER_89_631 VDD VSS sg13g2_decap_8
XFILLER_104_964 VDD VSS sg13g2_decap_8
XFILLER_89_664 VDD VSS sg13g2_decap_8
XFILLER_103_430 VDD VSS sg13g2_decap_8
XFILLER_107_63 VDD VSS sg13g2_decap_8
XFILLER_1_546 VDD VSS sg13g2_decap_8
XFILLER_77_837 VDD VSS sg13g2_decap_8
XFILLER_27_1057 VDD VSS sg13g2_decap_4
XFILLER_67_56 VDD VSS sg13g2_decap_8
XFILLER_103_496 VDD VSS sg13g2_decap_8
XFILLER_29_252 VDD VSS sg13g2_decap_8
XFILLER_18_959 VDD VSS sg13g2_decap_8
XFILLER_44_200 VDD VSS sg13g2_decap_8
XFILLER_83_77 VDD VSS sg13g2_decap_8
XFILLER_17_469 VDD VSS sg13g2_decap_8
XFILLER_32_406 VDD VSS sg13g2_decap_8
XFILLER_60_748 VDD VSS sg13g2_decap_8
XFILLER_73_1044 VDD VSS sg13g2_decap_8
XFILLER_41_951 VDD VSS sg13g2_decap_8
XFILLER_9_602 VDD VSS sg13g2_decap_8
XFILLER_8_112 VDD VSS sg13g2_decap_8
XFILLER_13_686 VDD VSS sg13g2_decap_8
XFILLER_40_461 VDD VSS sg13g2_decap_8
XFILLER_40_472 VDD VSS sg13g2_fill_1
XFILLER_12_196 VDD VSS sg13g2_decap_8
XFILLER_9_679 VDD VSS sg13g2_decap_8
XFILLER_32_70 VDD VSS sg13g2_decap_8
XFILLER_8_189 VDD VSS sg13g2_decap_8
XFILLER_10_1050 VDD VSS sg13g2_decap_8
XFILLER_59_7 VDD VSS sg13g2_decap_8
XFILLER_99_428 VDD VSS sg13g2_decap_8
X_1460_ VSS VDD _1382_/Y _1463_/B _2249_/D _1459_/Y sg13g2_a21oi_1
XFILLER_5_896 VDD VSS sg13g2_decap_8
X_1391_ _2267_/Q _1492_/A _2265_/Q _1409_/C _1391_/Y VDD VSS sg13g2_nor4_1
XFILLER_95_623 VDD VSS sg13g2_decap_8
XFILLER_68_848 VDD VSS sg13g2_decap_8
XFILLER_110_956 VDD VSS sg13g2_decap_8
XFILLER_79_196 VDD VSS sg13g2_decap_8
XFILLER_94_133 VDD VSS sg13g2_decap_8
XFILLER_67_336 VDD VSS sg13g2_decap_4
XFILLER_83_829 VDD VSS sg13g2_decap_8
XFILLER_82_306 VDD VSS sg13g2_decap_8
XFILLER_48_561 VDD VSS sg13g2_decap_8
X_2012_ _2011_/Y VDD _2321_/D VSS _2033_/B _2025_/A sg13g2_o21ai_1
XFILLER_82_328 VDD VSS sg13g2_decap_8
XFILLER_63_531 VDD VSS sg13g2_decap_8
XFILLER_36_756 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_51_737 VDD VSS sg13g2_decap_8
XFILLER_23_406 VDD VSS sg13g2_decap_8
XFILLER_35_266 VDD VSS sg13g2_decap_8
XFILLER_85_0 VDD VSS sg13g2_decap_8
XFILLER_32_973 VDD VSS sg13g2_decap_8
XFILLER_31_483 VDD VSS sg13g2_decap_8
XFILLER_105_728 VDD VSS sg13g2_decap_8
X_1727_ _1727_/Y _2230_/Q _2238_/Q VDD VSS sg13g2_nand2b_1
X_1658_ _1671_/C _1658_/B _2302_/D VDD VSS sg13g2_nor2_1
XFILLER_104_238 VDD VSS sg13g2_decap_8
XFILLER_86_623 VDD VSS sg13g2_decap_8
XFILLER_98_483 VDD VSS sg13g2_decap_8
XFILLER_59_826 VDD VSS sg13g2_fill_1
X_1589_ _1592_/B _1589_/A _1589_/B _1589_/C VDD VSS sg13g2_and3_1
XFILLER_101_956 VDD VSS sg13g2_decap_8
XFILLER_74_807 VDD VSS sg13g2_decap_8
XFILLER_85_122 VDD VSS sg13g2_fill_2
XFILLER_58_358 VDD VSS sg13g2_decap_8
XFILLER_100_455 VDD VSS sg13g2_decap_8
XFILLER_85_199 VDD VSS sg13g2_decap_8
XFILLER_2_1015 VDD VSS sg13g2_decap_8
XFILLER_57_1017 VDD VSS sg13g2_decap_8
XFILLER_27_756 VDD VSS sg13g2_decap_8
XFILLER_81_361 VDD VSS sg13g2_decap_8
XFILLER_14_406 VDD VSS sg13g2_decap_8
XFILLER_53_14 VDD VSS sg13g2_decap_4
XFILLER_26_266 VDD VSS sg13g2_decap_8
XFILLER_53_69 VDD VSS sg13g2_decap_8
XFILLER_23_973 VDD VSS sg13g2_decap_8
XFILLER_50_770 VDD VSS sg13g2_decap_8
XFILLER_10_623 VDD VSS sg13g2_decap_8
XFILLER_22_483 VDD VSS sg13g2_decap_8
XFILLER_33_1050 VDD VSS sg13g2_decap_8
XFILLER_6_616 VDD VSS sg13g2_decap_8
XFILLER_5_126 VDD VSS sg13g2_decap_8
XFILLER_108_577 VDD VSS sg13g2_decap_8
XFILLER_2_833 VDD VSS sg13g2_decap_8
XFILLER_104_750 VDD VSS sg13g2_decap_8
XFILLER_1_343 VDD VSS sg13g2_decap_8
XFILLER_78_77 VDD VSS sg13g2_decap_8
XFILLER_89_494 VDD VSS sg13g2_decap_8
XFILLER_76_133 VDD VSS sg13g2_decap_8
XFILLER_77_667 VDD VSS sg13g2_decap_8
XFILLER_94_21 VDD VSS sg13g2_decap_8
XFILLER_40_1054 VDD VSS sg13g2_decap_8
XFILLER_64_328 VDD VSS sg13g2_decap_8
XFILLER_64_339 VDD VSS sg13g2_fill_1
XFILLER_94_98 VDD VSS sg13g2_decap_8
XFILLER_45_553 VDD VSS sg13g2_decap_8
XFILLER_18_756 VDD VSS sg13g2_decap_8
XFILLER_27_70 VDD VSS sg13g2_decap_8
XFILLER_17_266 VDD VSS sg13g2_decap_8
XFILLER_32_203 VDD VSS sg13g2_decap_8
XFILLER_60_545 VDD VSS sg13g2_decap_8
XFILLER_14_973 VDD VSS sg13g2_decap_8
XFILLER_13_483 VDD VSS sg13g2_decap_8
XFILLER_43_91 VDD VSS sg13g2_decap_8
XFILLER_9_476 VDD VSS sg13g2_decap_8
X_1512_ VSS VDD _1510_/A _1510_/B _1513_/C hold530/X sg13g2_a21oi_1
XFILLER_5_693 VDD VSS sg13g2_decap_8
X_1443_ VDD _2241_/D _1443_/A VSS sg13g2_inv_1
XFILLER_87_409 VDD VSS sg13g2_decap_8
XFILLER_68_601 VDD VSS sg13g2_decap_8
XFILLER_4_63 VDD VSS sg13g2_decap_8
XFILLER_96_954 VDD VSS sg13g2_decap_8
XFILLER_95_420 VDD VSS sg13g2_decap_8
X_1374_ _1374_/Y _1374_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_68_645 VDD VSS sg13g2_decap_8
XFILLER_110_753 VDD VSS sg13g2_decap_8
XFILLER_83_626 VDD VSS sg13g2_decap_8
XFILLER_67_188 VDD VSS sg13g2_decap_8
XFILLER_64_851 VDD VSS sg13g2_decap_8
XFILLER_64_862 VDD VSS sg13g2_fill_1
XFILLER_36_553 VDD VSS sg13g2_decap_8
XFILLER_64_873 VDD VSS sg13g2_decap_8
XFILLER_51_523 VDD VSS sg13g2_decap_8
XFILLER_23_203 VDD VSS sg13g2_decap_8
XFILLER_63_394 VDD VSS sg13g2_decap_8
XFILLER_56_1050 VDD VSS sg13g2_decap_8
XFILLER_32_770 VDD VSS sg13g2_decap_8
XFILLER_20_910 VDD VSS sg13g2_decap_8
XFILLER_17_1001 VDD VSS sg13g2_decap_8
XFILLER_23_28 VDD VSS sg13g2_decap_8
XFILLER_31_280 VDD VSS sg13g2_decap_8
XFILLER_104_1048 VDD VSS sg13g2_decap_8
XFILLER_104_1059 VDD VSS sg13g2_fill_2
XFILLER_20_987 VDD VSS sg13g2_decap_8
XFILLER_105_547 VDD VSS sg13g2_fill_1
XFILLER_87_910 VDD VSS sg13g2_decap_8
XFILLER_63_1010 VDD VSS sg13g2_decap_4
XFILLER_59_623 VDD VSS sg13g2_decap_8
XFILLER_48_14 VDD VSS sg13g2_decap_8
XFILLER_58_100 VDD VSS sg13g2_decap_8
XFILLER_111_1008 VDD VSS sg13g2_decap_8
XFILLER_86_475 VDD VSS sg13g2_decap_8
XFILLER_59_678 VDD VSS sg13g2_decap_8
XFILLER_101_786 VDD VSS sg13g2_decap_8
XFILLER_104_42 VDD VSS sg13g2_decap_8
XFILLER_39_380 VDD VSS sg13g2_decap_8
XFILLER_73_136 VDD VSS sg13g2_decap_8
XFILLER_27_553 VDD VSS sg13g2_decap_8
XFILLER_64_35 VDD VSS sg13g2_decap_8
XFILLER_82_681 VDD VSS sg13g2_decap_8
X_2218__104 VDD VSS _2218_/RESET_B sg13g2_tiehi
XFILLER_55_895 VDD VSS sg13g2_decap_8
XFILLER_14_203 VDD VSS sg13g2_decap_8
XFILLER_70_843 VDD VSS sg13g2_decap_8
Xfanout40 _1264_/X fanout40/X VDD VSS sg13g2_buf_1
XFILLER_30_707 VDD VSS sg13g2_decap_8
XFILLER_11_910 VDD VSS sg13g2_decap_8
XFILLER_80_56 VDD VSS sg13g2_decap_8
Xfanout62 _2124_/A _2144_/S0 VDD VSS sg13g2_buf_1
XFILLER_23_770 VDD VSS sg13g2_decap_8
XFILLER_10_420 VDD VSS sg13g2_decap_8
Xfanout73 _2107_/B1 _1236_/C VDD VSS sg13g2_buf_1
Xfanout51 _2287_/Q _1589_/B VDD VSS sg13g2_buf_1
XFILLER_70_1058 VDD VSS sg13g2_fill_2
XFILLER_7_903 VDD VSS sg13g2_decap_8
XFILLER_22_280 VDD VSS sg13g2_decap_8
XFILLER_6_413 VDD VSS sg13g2_decap_8
XFILLER_11_987 VDD VSS sg13g2_decap_8
XFILLER_109_875 VDD VSS sg13g2_decap_8
XFILLER_89_21 VDD VSS sg13g2_decap_8
XFILLER_10_497 VDD VSS sg13g2_decap_8
XFILLER_89_98 VDD VSS sg13g2_decap_8
XFILLER_2_630 VDD VSS sg13g2_decap_8
XFILLER_97_729 VDD VSS sg13g2_decap_4
XFILLER_96_217 VDD VSS sg13g2_decap_8
XFILLER_1_140 VDD VSS sg13g2_decap_8
XFILLER_78_965 VDD VSS sg13g2_decap_8
XFILLER_104_591 VDD VSS sg13g2_decap_8
XFILLER_111_539 VDD VSS sg13g2_decap_8
XFILLER_77_475 VDD VSS sg13g2_decap_8
XFILLER_38_807 VDD VSS sg13g2_decap_8
XFILLER_49_133 VDD VSS sg13g2_decap_8
XFILLER_92_434 VDD VSS sg13g2_decap_8
XFILLER_93_979 VDD VSS sg13g2_fill_2
XFILLER_18_553 VDD VSS sg13g2_decap_8
XFILLER_38_91 VDD VSS sg13g2_decap_8
XFILLER_64_136 VDD VSS sg13g2_decap_8
XFILLER_46_873 VDD VSS sg13g2_decap_8
XFILLER_45_350 VDD VSS sg13g2_decap_4
XFILLER_60_331 VDD VSS sg13g2_decap_8
XFILLER_61_865 VDD VSS sg13g2_decap_8
XFILLER_33_567 VDD VSS sg13g2_decap_8
XFILLER_21_707 VDD VSS sg13g2_decap_8
X_1992_ _2005_/C _1992_/A _1992_/B VDD VSS sg13g2_xnor2_1
XFILLER_60_375 VDD VSS sg13g2_decap_8
XFILLER_20_217 VDD VSS sg13g2_decap_8
XFILLER_14_770 VDD VSS sg13g2_decap_8
XFILLER_13_280 VDD VSS sg13g2_decap_8
Xclkload10 clkload10/Y _2373_/CLK VDD VSS sg13g2_inv_2
XFILLER_9_273 VDD VSS sg13g2_decap_8
XFILLER_6_980 VDD VSS sg13g2_decap_8
XFILLER_88_707 VDD VSS sg13g2_decap_8
XFILLER_47_1027 VDD VSS sg13g2_decap_8
XFILLER_5_490 VDD VSS sg13g2_decap_8
XFILLER_48_0 VDD VSS sg13g2_decap_8
XFILLER_88_729 VDD VSS sg13g2_decap_8
XFILLER_102_528 VDD VSS sg13g2_decap_8
XFILLER_69_943 VDD VSS sg13g2_decap_8
X_1426_ _1426_/Y _1426_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_68_420 VDD VSS sg13g2_decap_8
XFILLER_110_550 VDD VSS sg13g2_decap_8
XFILLER_84_913 VDD VSS sg13g2_decap_4
X_1357_ VDD _2207_/D _1357_/A VSS sg13g2_inv_1
XFILLER_95_272 VDD VSS sg13g2_decap_8
XFILLER_56_637 VDD VSS sg13g2_decap_8
XFILLER_18_28 VDD VSS sg13g2_decap_8
X_1288_ _1288_/Y _1322_/B1 hold355/X _1322_/A2 _2338_/Q VDD VSS sg13g2_a22oi_1
XFILLER_83_445 VDD VSS sg13g2_decap_8
XFILLER_37_840 VDD VSS sg13g2_decap_8
XFILLER_55_147 VDD VSS sg13g2_decap_8
XFILLER_52_810 VDD VSS sg13g2_decap_8
XFILLER_36_350 VDD VSS sg13g2_decap_8
XFILLER_24_567 VDD VSS sg13g2_decap_8
XFILLER_12_707 VDD VSS sg13g2_decap_8
XFILLER_34_49 VDD VSS sg13g2_decap_8
XFILLER_11_217 VDD VSS sg13g2_decap_8
XFILLER_109_105 VDD VSS sg13g2_decap_8
Xclkload4 VDD clkload4/Y clkload4/A VSS sg13g2_inv_1
XFILLER_20_784 VDD VSS sg13g2_decap_8
XFILLER_4_917 VDD VSS sg13g2_decap_8
XFILLER_3_427 VDD VSS sg13g2_decap_8
XFILLER_106_867 VDD VSS sg13g2_decap_8
XFILLER_105_344 VDD VSS sg13g2_decap_8
XFILLER_79_729 VDD VSS sg13g2_decap_8
XFILLER_78_206 VDD VSS sg13g2_fill_1
XFILLER_59_57 VDD VSS sg13g2_fill_2
XFILLER_59_68 VDD VSS sg13g2_decap_8
XFILLER_78_239 VDD VSS sg13g2_decap_8
XFILLER_87_773 VDD VSS sg13g2_decap_8
XFILLER_8_1043 VDD VSS sg13g2_decap_8
XFILLER_101_594 VDD VSS sg13g2_decap_8
XFILLER_101_561 VDD VSS sg13g2_fill_1
XFILLER_47_637 VDD VSS sg13g2_decap_8
XFILLER_59_497 VDD VSS sg13g2_decap_8
XFILLER_90_916 VDD VSS sg13g2_decap_8
XFILLER_75_56 VDD VSS sg13g2_decap_8
XFILLER_28_840 VDD VSS sg13g2_decap_8
XFILLER_43_821 VDD VSS sg13g2_decap_8
XFILLER_27_350 VDD VSS sg13g2_decap_8
XFILLER_70_640 VDD VSS sg13g2_decap_8
XFILLER_55_692 VDD VSS sg13g2_decap_8
XFILLER_15_567 VDD VSS sg13g2_decap_8
XFILLER_30_504 VDD VSS sg13g2_decap_8
XFILLER_91_77 VDD VSS sg13g2_decap_8
XFILLER_43_898 VDD VSS sg13g2_decap_8
XFILLER_7_700 VDD VSS sg13g2_decap_8
XFILLER_6_210 VDD VSS sg13g2_decap_8
XFILLER_11_784 VDD VSS sg13g2_decap_8
XFILLER_10_294 VDD VSS sg13g2_decap_8
XFILLER_7_777 VDD VSS sg13g2_decap_8
XFILLER_109_672 VDD VSS sg13g2_decap_8
XFILLER_6_287 VDD VSS sg13g2_decap_8
XFILLER_40_70 VDD VSS sg13g2_decap_8
XFILLER_112_826 VDD VSS sg13g2_decap_8
XFILLER_41_7 VDD VSS sg13g2_decap_8
XFILLER_111_336 VDD VSS sg13g2_decap_8
X_2260_ _2260_/RESET_B VSS VDD _2260_/D _2260_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_3_994 VDD VSS sg13g2_decap_8
XFILLER_38_604 VDD VSS sg13g2_decap_8
X_1211_ VDD _1211_/Y _2248_/Q VSS sg13g2_inv_1
X_2191_ _2191_/RESET_B VSS VDD _2191_/D _2191_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_93_710 VDD VSS sg13g2_decap_8
XFILLER_66_935 VDD VSS sg13g2_decap_8
XFILLER_92_242 VDD VSS sg13g2_decap_8
XFILLER_77_294 VDD VSS sg13g2_decap_8
XFILLER_65_445 VDD VSS sg13g2_decap_8
XFILLER_1_42 VDD VSS sg13g2_decap_8
XFILLER_19_840 VDD VSS sg13g2_decap_8
XFILLER_37_147 VDD VSS sg13g2_decap_8
XFILLER_93_787 VDD VSS sg13g2_decap_8
XFILLER_93_798 VDD VSS sg13g2_fill_2
XFILLER_80_404 VDD VSS sg13g2_decap_8
XFILLER_18_350 VDD VSS sg13g2_decap_8
XFILLER_92_286 VDD VSS sg13g2_fill_1
XFILLER_34_854 VDD VSS sg13g2_decap_8
XFILLER_52_117 VDD VSS sg13g2_decap_8
XFILLER_21_504 VDD VSS sg13g2_decap_8
XFILLER_33_364 VDD VSS sg13g2_decap_8
XFILLER_61_695 VDD VSS sg13g2_fill_2
XFILLER_60_161 VDD VSS sg13g2_decap_4
X_1975_ _1975_/Y _1976_/A _1976_/B VDD VSS sg13g2_nand2_1
XFILLER_14_1015 VDD VSS sg13g2_decap_8
XFILLER_106_119 VDD VSS sg13g2_decap_8
XFILLER_102_303 VDD VSS sg13g2_fill_1
XFILLER_88_537 VDD VSS sg13g2_decap_4
XFILLER_69_762 VDD VSS sg13g2_decap_8
X_1409_ _2267_/Q _2266_/Q _1409_/C _1410_/B VDD VSS sg13g2_nor3_1
XFILLER_29_49 VDD VSS sg13g2_decap_8
XFILLER_96_592 VDD VSS sg13g2_decap_8
XFILLER_60_1046 VDD VSS sg13g2_decap_8
XFILLER_21_1008 VDD VSS sg13g2_decap_8
XFILLER_29_637 VDD VSS sg13g2_decap_8
XFILLER_56_412 VDD VSS sg13g2_decap_8
XFILLER_72_905 VDD VSS sg13g2_decap_8
XFILLER_83_231 VDD VSS sg13g2_decap_8
XFILLER_83_220 VDD VSS sg13g2_fill_2
XFILLER_57_979 VDD VSS sg13g2_decap_8
XFILLER_28_147 VDD VSS sg13g2_decap_8
XFILLER_72_916 VDD VSS sg13g2_fill_2
XFILLER_71_404 VDD VSS sg13g2_decap_8
XFILLER_101_21 VDD VSS sg13g2_decap_8
XFILLER_40_802 VDD VSS sg13g2_decap_8
XFILLER_25_854 VDD VSS sg13g2_decap_8
XFILLER_52_684 VDD VSS sg13g2_decap_8
XFILLER_12_504 VDD VSS sg13g2_decap_8
XFILLER_51_150 VDD VSS sg13g2_decap_8
XFILLER_61_14 VDD VSS sg13g2_decap_8
XFILLER_24_364 VDD VSS sg13g2_decap_8
XFILLER_101_98 VDD VSS sg13g2_decap_8
XFILLER_40_879 VDD VSS sg13g2_decap_8
XFILLER_20_581 VDD VSS sg13g2_decap_8
XFILLER_4_714 VDD VSS sg13g2_decap_8
XFILLER_3_224 VDD VSS sg13g2_decap_8
XFILLER_106_664 VDD VSS sg13g2_decap_8
XFILLER_105_185 VDD VSS sg13g2_fill_2
XFILLER_79_526 VDD VSS sg13g2_decap_8
XFILLER_10_84 VDD VSS sg13g2_decap_8
XFILLER_0_931 VDD VSS sg13g2_decap_8
XFILLER_66_209 VDD VSS sg13g2_decap_8
XFILLER_102_881 VDD VSS sg13g2_decap_8
XFILLER_75_721 VDD VSS sg13g2_decap_8
XFILLER_94_529 VDD VSS sg13g2_decap_8
XFILLER_86_77 VDD VSS sg13g2_decap_8
XFILLER_59_250 VDD VSS sg13g2_fill_2
XFILLER_59_272 VDD VSS sg13g2_fill_2
XFILLER_19_147 VDD VSS sg13g2_decap_8
XFILLER_90_724 VDD VSS sg13g2_decap_8
XFILLER_47_467 VDD VSS sg13g2_fill_1
XFILLER_74_286 VDD VSS sg13g2_decap_8
XFILLER_63_949 VDD VSS sg13g2_decap_8
XFILLER_37_1015 VDD VSS sg13g2_decap_8
XFILLER_16_854 VDD VSS sg13g2_decap_8
XFILLER_35_70 VDD VSS sg13g2_decap_8
XFILLER_70_470 VDD VSS sg13g2_decap_8
XFILLER_43_695 VDD VSS sg13g2_decap_8
XFILLER_15_364 VDD VSS sg13g2_decap_8
XFILLER_30_301 VDD VSS sg13g2_decap_8
XFILLER_89_7 VDD VSS sg13g2_decap_8
XFILLER_31_868 VDD VSS sg13g2_decap_8
X_1760_ _1770_/A _1760_/A _1760_/B VDD VSS sg13g2_nand2_1
XFILLER_30_378 VDD VSS sg13g2_decap_8
XFILLER_11_581 VDD VSS sg13g2_decap_8
X_1691_ _1692_/B _2314_/Q _2300_/Q VDD VSS sg13g2_xnor2_1
Xhold508 _2267_/Q VDD VSS _1495_/A sg13g2_dlygate4sd3_1
XFILLER_7_574 VDD VSS sg13g2_decap_8
Xhold519 _2244_/Q VDD VSS _1449_/A sg13g2_dlygate4sd3_1
XFILLER_83_1024 VDD VSS sg13g2_decap_8
XFILLER_98_813 VDD VSS sg13g2_decap_8
XFILLER_97_301 VDD VSS sg13g2_decap_8
XFILLER_112_623 VDD VSS sg13g2_decap_8
XFILLER_44_1019 VDD VSS sg13g2_decap_8
X_2312_ _2312_/RESET_B VSS VDD _2312_/D _2312_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_3_791 VDD VSS sg13g2_decap_8
XFILLER_111_133 VDD VSS sg13g2_decap_8
X_2243_ _2243_/RESET_B VSS VDD _2243_/D _2243_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_39_913 VDD VSS sg13g2_decap_8
X_2174_ _2174_/RESET_B VSS VDD _2174_/D _2174_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_78_592 VDD VSS sg13g2_decap_4
XFILLER_54_927 VDD VSS sg13g2_decap_8
XFILLER_38_467 VDD VSS sg13g2_decap_8
XFILLER_80_234 VDD VSS sg13g2_decap_8
XFILLER_62_960 VDD VSS sg13g2_decap_8
XFILLER_34_651 VDD VSS sg13g2_decap_8
XFILLER_61_481 VDD VSS sg13g2_decap_8
XFILLER_33_161 VDD VSS sg13g2_decap_8
XFILLER_21_301 VDD VSS sg13g2_decap_8
XFILLER_22_868 VDD VSS sg13g2_decap_8
XFILLER_21_378 VDD VSS sg13g2_decap_8
X_1958_ _1978_/C _1958_/A _1958_/B VDD VSS sg13g2_xnor2_1
XFILLER_31_28 VDD VSS sg13g2_decap_8
X_1889_ _1891_/B _1889_/A _1889_/B VDD VSS sg13g2_xnor2_1
XFILLER_89_824 VDD VSS sg13g2_decap_4
XFILLER_103_623 VDD VSS sg13g2_decap_8
XFILLER_88_312 VDD VSS sg13g2_decap_4
XFILLER_1_728 VDD VSS sg13g2_decap_8
XFILLER_102_133 VDD VSS sg13g2_decap_8
XFILLER_0_238 VDD VSS sg13g2_decap_8
XFILLER_56_14 VDD VSS sg13g2_decap_8
XFILLER_99_1031 VDD VSS sg13g2_decap_8
XFILLER_5_1057 VDD VSS sg13g2_decap_4
XFILLER_29_434 VDD VSS sg13g2_decap_8
XFILLER_57_765 VDD VSS sg13g2_decap_8
XFILLER_56_242 VDD VSS sg13g2_decap_8
XFILLER_56_58 VDD VSS sg13g2_decap_4
XFILLER_72_724 VDD VSS sg13g2_fill_2
XFILLER_71_212 VDD VSS sg13g2_decap_8
XFILLER_112_42 VDD VSS sg13g2_decap_8
XFILLER_71_256 VDD VSS sg13g2_decap_8
XFILLER_25_651 VDD VSS sg13g2_decap_8
XFILLER_72_35 VDD VSS sg13g2_decap_8
XFILLER_12_301 VDD VSS sg13g2_decap_8
XFILLER_24_161 VDD VSS sg13g2_decap_8
XFILLER_52_481 VDD VSS sg13g2_decap_8
XFILLER_13_868 VDD VSS sg13g2_decap_8
XFILLER_40_676 VDD VSS sg13g2_decap_8
XFILLER_12_378 VDD VSS sg13g2_decap_8
XFILLER_107_940 VDD VSS sg13g2_decap_8
XFILLER_4_511 VDD VSS sg13g2_decap_8
XFILLER_97_21 VDD VSS sg13g2_decap_8
XFILLER_4_588 VDD VSS sg13g2_decap_8
XFILLER_79_334 VDD VSS sg13g2_decap_8
XFILLER_97_98 VDD VSS sg13g2_decap_8
XFILLER_67_518 VDD VSS sg13g2_decap_8
XFILLER_94_359 VDD VSS sg13g2_decap_4
XFILLER_43_1052 VDD VSS sg13g2_decap_8
XFILLER_48_754 VDD VSS sg13g2_decap_8
XFILLER_47_231 VDD VSS sg13g2_decap_8
XFILLER_36_938 VDD VSS sg13g2_decap_8
XFILLER_47_264 VDD VSS sg13g2_decap_8
XFILLER_75_595 VDD VSS sg13g2_decap_8
XFILLER_63_779 VDD VSS sg13g2_decap_8
XFILLER_62_234 VDD VSS sg13g2_fill_2
XFILLER_16_651 VDD VSS sg13g2_decap_8
XFILLER_46_91 VDD VSS sg13g2_decap_8
XFILLER_35_448 VDD VSS sg13g2_decap_8
XFILLER_90_587 VDD VSS sg13g2_decap_8
XFILLER_15_161 VDD VSS sg13g2_decap_8
XFILLER_31_665 VDD VSS sg13g2_decap_8
X_1812_ _1812_/B _1812_/A _1949_/A VDD VSS sg13g2_xor2_1
XFILLER_50_1045 VDD VSS sg13g2_decap_8
XFILLER_30_175 VDD VSS sg13g2_decap_8
X_1743_ _1774_/A _1772_/A _1750_/A VDD VSS sg13g2_nor2_1
XFILLER_7_63 VDD VSS sg13g2_decap_8
XFILLER_8_861 VDD VSS sg13g2_decap_8
XFILLER_11_1029 VDD VSS sg13g2_decap_8
Xhold305 _1322_/Y VDD VSS _1323_/A sg13g2_dlygate4sd3_1
Xhold316 _2201_/Q VDD VSS hold316/X sg13g2_dlygate4sd3_1
X_1674_ _1674_/A _1674_/B _1677_/B VDD VSS sg13g2_and2_1
XFILLER_7_371 VDD VSS sg13g2_decap_8
Xhold327 _2186_/Q VDD VSS hold327/X sg13g2_dlygate4sd3_1
Xhold338 _2187_/Q VDD VSS hold338/X sg13g2_dlygate4sd3_1
Xhold349 _2256_/Q VDD VSS _1242_/B sg13g2_dlygate4sd3_1
X_2283__171 VDD VSS _2283_/RESET_B sg13g2_tiehi
XFILLER_86_816 VDD VSS sg13g2_decap_8
XFILLER_112_420 VDD VSS sg13g2_decap_8
XFILLER_30_0 VDD VSS sg13g2_decap_8
XFILLER_97_186 VDD VSS sg13g2_decap_8
XFILLER_39_710 VDD VSS sg13g2_decap_8
XFILLER_58_518 VDD VSS sg13g2_decap_8
XFILLER_100_637 VDD VSS sg13g2_decap_8
XFILLER_112_497 VDD VSS sg13g2_decap_8
X_2226_ _2226__88/L_HI VSS VDD _2226_/D _2226_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_85_348 VDD VSS sg13g2_decap_8
XFILLER_94_871 VDD VSS sg13g2_decap_8
XFILLER_39_787 VDD VSS sg13g2_decap_8
XFILLER_66_540 VDD VSS sg13g2_decap_8
XFILLER_38_231 VDD VSS sg13g2_decap_8
X_2157_ _2162_/A _2162_/B _2345_/D VDD VSS sg13g2_nor2_1
XFILLER_81_510 VDD VSS sg13g2_decap_8
XFILLER_27_938 VDD VSS sg13g2_decap_8
XFILLER_54_735 VDD VSS sg13g2_fill_1
XFILLER_26_28 VDD VSS sg13g2_decap_8
X_2088_ _2086_/Y VDD _2342_/D VSS _2156_/A _2087_/Y sg13g2_o21ai_1
XFILLER_53_245 VDD VSS sg13g2_decap_8
XFILLER_26_448 VDD VSS sg13g2_decap_8
XFILLER_81_587 VDD VSS sg13g2_decap_8
XFILLER_107_1024 VDD VSS sg13g2_decap_8
XFILLER_50_974 VDD VSS sg13g2_decap_8
XFILLER_22_665 VDD VSS sg13g2_decap_8
XFILLER_10_805 VDD VSS sg13g2_decap_8
XFILLER_42_49 VDD VSS sg13g2_decap_8
XFILLER_21_175 VDD VSS sg13g2_decap_8
XFILLER_5_308 VDD VSS sg13g2_decap_8
XFILLER_108_759 VDD VSS sg13g2_decap_8
XFILLER_1_525 VDD VSS sg13g2_decap_8
XFILLER_104_943 VDD VSS sg13g2_decap_8
XFILLER_107_42 VDD VSS sg13g2_decap_8
XFILLER_27_1036 VDD VSS sg13g2_decap_8
XFILLER_77_816 VDD VSS sg13g2_decap_8
XFILLER_103_475 VDD VSS sg13g2_decap_8
XFILLER_67_35 VDD VSS sg13g2_decap_8
XFILLER_49_507 VDD VSS sg13g2_decap_8
XFILLER_76_359 VDD VSS sg13g2_fill_1
XFILLER_92_819 VDD VSS sg13g2_decap_8
XFILLER_57_551 VDD VSS sg13g2_decap_8
XFILLER_29_231 VDD VSS sg13g2_decap_8
XFILLER_18_938 VDD VSS sg13g2_decap_8
XFILLER_72_543 VDD VSS sg13g2_decap_8
XFILLER_84_392 VDD VSS sg13g2_decap_8
XFILLER_83_56 VDD VSS sg13g2_decap_8
XFILLER_17_448 VDD VSS sg13g2_decap_8
XFILLER_44_234 VDD VSS sg13g2_fill_1
XFILLER_72_598 VDD VSS sg13g2_decap_8
XFILLER_73_1023 VDD VSS sg13g2_decap_8
XFILLER_41_930 VDD VSS sg13g2_decap_8
XFILLER_34_1029 VDD VSS sg13g2_decap_8
XFILLER_13_665 VDD VSS sg13g2_decap_8
XFILLER_40_440 VDD VSS sg13g2_decap_8
XFILLER_12_175 VDD VSS sg13g2_decap_8
XFILLER_9_658 VDD VSS sg13g2_decap_8
XFILLER_40_484 VDD VSS sg13g2_decap_8
XFILLER_8_168 VDD VSS sg13g2_decap_8
XFILLER_5_875 VDD VSS sg13g2_decap_8
XFILLER_4_385 VDD VSS sg13g2_decap_8
XFILLER_106_280 VDD VSS sg13g2_fill_1
X_1390_ _1389_/Y VDD _1390_/Y VSS _1366_/Y _1388_/Y sg13g2_o21ai_1
XFILLER_110_935 VDD VSS sg13g2_decap_8
XFILLER_68_827 VDD VSS sg13g2_decap_8
XFILLER_67_315 VDD VSS sg13g2_decap_8
XFILLER_83_808 VDD VSS sg13g2_decap_8
XFILLER_94_112 VDD VSS sg13g2_decap_8
XFILLER_95_679 VDD VSS sg13g2_decap_8
X_2011_ _2011_/Y _2074_/A _2031_/A VDD VSS sg13g2_nand2_1
XFILLER_76_893 VDD VSS sg13g2_decap_8
XFILLER_94_189 VDD VSS sg13g2_decap_8
XFILLER_36_735 VDD VSS sg13g2_decap_8
XFILLER_63_510 VDD VSS sg13g2_decap_8
XFILLER_90_340 VDD VSS sg13g2_decap_8
XFILLER_35_245 VDD VSS sg13g2_decap_8
XFILLER_32_952 VDD VSS sg13g2_decap_8
XFILLER_31_462 VDD VSS sg13g2_decap_8
XFILLER_50_259 VDD VSS sg13g2_decap_8
XFILLER_78_0 VDD VSS sg13g2_decap_8
XFILLER_105_707 VDD VSS sg13g2_decap_8
X_1726_ _1760_/A _1726_/A _2242_/Q VDD VSS sg13g2_nand2_1
X_1657_ _1657_/Y _1646_/Y _1656_/X hold435/X _1671_/B VDD VSS sg13g2_a22oi_1
XFILLER_104_217 VDD VSS sg13g2_decap_8
XFILLER_99_952 VDD VSS sg13g2_fill_2
X_1588_ VSS VDD _1589_/A _1589_/C _1590_/B _1589_/B sg13g2_a21oi_1
XFILLER_98_462 VDD VSS sg13g2_decap_8
XFILLER_101_935 VDD VSS sg13g2_decap_8
XFILLER_112_294 VDD VSS sg13g2_decap_8
XFILLER_100_412 VDD VSS sg13g2_fill_1
XFILLER_58_337 VDD VSS sg13g2_decap_8
XFILLER_86_679 VDD VSS sg13g2_decap_8
XFILLER_37_49 VDD VSS sg13g2_decap_8
XFILLER_85_178 VDD VSS sg13g2_decap_8
XFILLER_39_584 VDD VSS sg13g2_decap_8
XFILLER_27_735 VDD VSS sg13g2_decap_8
X_2209_ _2209_/RESET_B VSS VDD _2209_/D _2209_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_82_841 VDD VSS sg13g2_decap_8
XFILLER_81_340 VDD VSS sg13g2_decap_8
X_2179__182 VDD VSS _2179_/RESET_B sg13g2_tiehi
XFILLER_66_392 VDD VSS sg13g2_decap_8
XFILLER_54_532 VDD VSS sg13g2_decap_4
XFILLER_26_245 VDD VSS sg13g2_decap_8
XFILLER_23_952 VDD VSS sg13g2_decap_8
XFILLER_42_749 VDD VSS sg13g2_decap_8
XFILLER_41_226 VDD VSS sg13g2_decap_4
XFILLER_41_248 VDD VSS sg13g2_decap_8
XFILLER_10_602 VDD VSS sg13g2_decap_8
XFILLER_22_462 VDD VSS sg13g2_decap_8
XFILLER_108_501 VDD VSS sg13g2_decap_8
XFILLER_5_105 VDD VSS sg13g2_decap_8
XFILLER_10_679 VDD VSS sg13g2_decap_8
XFILLER_108_556 VDD VSS sg13g2_decap_8
XFILLER_2_812 VDD VSS sg13g2_decap_8
XFILLER_78_56 VDD VSS sg13g2_decap_8
XFILLER_1_322 VDD VSS sg13g2_decap_8
XFILLER_89_451 VDD VSS sg13g2_decap_8
XFILLER_89_462 VDD VSS sg13g2_decap_4
XFILLER_2_889 VDD VSS sg13g2_decap_8
XFILLER_77_646 VDD VSS sg13g2_decap_8
XFILLER_76_112 VDD VSS sg13g2_decap_8
XFILLER_1_399 VDD VSS sg13g2_decap_8
XFILLER_49_337 VDD VSS sg13g2_decap_8
XFILLER_64_307 VDD VSS sg13g2_decap_8
XFILLER_76_189 VDD VSS sg13g2_decap_8
XFILLER_94_77 VDD VSS sg13g2_decap_8
XFILLER_40_1033 VDD VSS sg13g2_decap_8
XFILLER_18_735 VDD VSS sg13g2_decap_8
XFILLER_17_245 VDD VSS sg13g2_decap_8
XFILLER_45_532 VDD VSS sg13g2_decap_8
XFILLER_72_373 VDD VSS sg13g2_decap_8
Xclkbuf_2_0__f_clk clkbuf_leaf_0_clk/A clkbuf_0_clk/X VDD VSS sg13g2_buf_16
XFILLER_33_749 VDD VSS sg13g2_decap_8
XFILLER_60_524 VDD VSS sg13g2_decap_8
XFILLER_14_952 VDD VSS sg13g2_decap_8
XFILLER_32_259 VDD VSS sg13g2_decap_8
XFILLER_13_462 VDD VSS sg13g2_decap_8
XFILLER_43_70 VDD VSS sg13g2_decap_8
XFILLER_71_7 VDD VSS sg13g2_decap_8
XFILLER_9_455 VDD VSS sg13g2_decap_8
X_1511_ _1513_/B _1507_/Y _1516_/B _1503_/X hold530/X VDD VSS sg13g2_a22oi_1
XFILLER_5_672 VDD VSS sg13g2_decap_8
X_1442_ _1443_/A _1429_/Y hold480/X _1429_/B _1385_/A VDD VSS sg13g2_a22oi_1
XFILLER_4_182 VDD VSS sg13g2_decap_8
XFILLER_4_42 VDD VSS sg13g2_decap_8
XFILLER_96_933 VDD VSS sg13g2_decap_8
XFILLER_110_732 VDD VSS sg13g2_decap_8
X_1373_ _1373_/Y _1373_/A _1465_/C VDD VSS sg13g2_nand2_1
XFILLER_67_112 VDD VSS sg13g2_decap_8
XFILLER_96_999 VDD VSS sg13g2_fill_2
XFILLER_83_605 VDD VSS sg13g2_decap_8
XFILLER_95_476 VDD VSS sg13g2_decap_8
XFILLER_67_167 VDD VSS sg13g2_decap_8
XFILLER_64_830 VDD VSS sg13g2_decap_8
XFILLER_55_329 VDD VSS sg13g2_decap_8
XFILLER_36_532 VDD VSS sg13g2_decap_8
XFILLER_48_381 VDD VSS sg13g2_decap_8
XFILLER_63_373 VDD VSS sg13g2_decap_8
XFILLER_90_181 VDD VSS sg13g2_decap_8
XFILLER_24_749 VDD VSS sg13g2_decap_8
XFILLER_51_579 VDD VSS sg13g2_decap_8
XFILLER_23_259 VDD VSS sg13g2_decap_8
XFILLER_17_1057 VDD VSS sg13g2_decap_4
XFILLER_104_1027 VDD VSS sg13g2_decap_8
XFILLER_20_966 VDD VSS sg13g2_decap_8
XFILLER_3_609 VDD VSS sg13g2_decap_8
X_1709_ _1710_/B _1709_/A _1714_/A VDD VSS sg13g2_xnor2_1
XFILLER_105_526 VDD VSS sg13g2_decap_8
XFILLER_2_119 VDD VSS sg13g2_decap_8
XFILLER_98_281 VDD VSS sg13g2_decap_4
XFILLER_63_1044 VDD VSS sg13g2_decap_8
XFILLER_101_765 VDD VSS sg13g2_decap_8
XFILLER_86_454 VDD VSS sg13g2_decap_8
XFILLER_104_21 VDD VSS sg13g2_decap_8
XFILLER_100_275 VDD VSS sg13g2_decap_8
XFILLER_100_286 VDD VSS sg13g2_fill_2
XFILLER_73_126 VDD VSS sg13g2_decap_4
XFILLER_64_14 VDD VSS sg13g2_decap_8
XFILLER_27_532 VDD VSS sg13g2_decap_8
XFILLER_82_660 VDD VSS sg13g2_decap_8
XFILLER_70_822 VDD VSS sg13g2_decap_8
XFILLER_104_98 VDD VSS sg13g2_decap_8
XFILLER_55_874 VDD VSS sg13g2_decap_8
XFILLER_54_373 VDD VSS sg13g2_decap_8
XFILLER_42_513 VDD VSS sg13g2_decap_8
XFILLER_81_181 VDD VSS sg13g2_decap_8
XFILLER_54_384 VDD VSS sg13g2_fill_1
XFILLER_15_749 VDD VSS sg13g2_decap_8
Xfanout30 _1366_/Y _1367_/B VDD VSS sg13g2_buf_1
XFILLER_14_259 VDD VSS sg13g2_decap_8
XFILLER_70_1004 VDD VSS sg13g2_decap_8
XFILLER_70_899 VDD VSS sg13g2_decap_8
XFILLER_80_35 VDD VSS sg13g2_decap_8
Xfanout41 _1206_/Y _2124_/B VDD VSS sg13g2_buf_1
Xfanout63 _2269_/Q _2124_/A VDD VSS sg13g2_buf_1
Xfanout52 _1580_/A1 _1573_/A1 VDD VSS sg13g2_buf_1
Xfanout74 fanout78/A _2107_/B1 VDD VSS sg13g2_buf_1
XFILLER_11_966 VDD VSS sg13g2_decap_8
XFILLER_10_476 VDD VSS sg13g2_decap_8
XFILLER_13_84 VDD VSS sg13g2_decap_8
XFILLER_7_959 VDD VSS sg13g2_decap_8
XFILLER_109_854 VDD VSS sg13g2_decap_8
XFILLER_6_469 VDD VSS sg13g2_decap_8
XFILLER_108_364 VDD VSS sg13g2_fill_2
XFILLER_89_77 VDD VSS sg13g2_decap_8
XFILLER_8_0 VDD VSS sg13g2_decap_8
XFILLER_111_518 VDD VSS sg13g2_decap_8
XFILLER_78_944 VDD VSS sg13g2_decap_8
XFILLER_104_570 VDD VSS sg13g2_decap_8
XFILLER_2_686 VDD VSS sg13g2_decap_8
XFILLER_77_443 VDD VSS sg13g2_fill_2
XFILLER_77_454 VDD VSS sg13g2_decap_8
XFILLER_65_605 VDD VSS sg13g2_fill_2
XFILLER_1_196 VDD VSS sg13g2_decap_8
XFILLER_93_958 VDD VSS sg13g2_decap_8
XFILLER_38_70 VDD VSS sg13g2_decap_8
XFILLER_37_329 VDD VSS sg13g2_decap_8
XFILLER_49_189 VDD VSS sg13g2_decap_8
XFILLER_18_532 VDD VSS sg13g2_decap_8
XFILLER_73_660 VDD VSS sg13g2_fill_1
XFILLER_61_811 VDD VSS sg13g2_decap_8
XFILLER_61_822 VDD VSS sg13g2_fill_1
XFILLER_73_693 VDD VSS sg13g2_decap_8
XFILLER_61_844 VDD VSS sg13g2_decap_8
XFILLER_33_546 VDD VSS sg13g2_decap_8
XFILLER_45_395 VDD VSS sg13g2_decap_8
X_1991_ _1971_/C _1971_/B _1971_/A _1991_/X VDD VSS sg13g2_a21o_1
XFILLER_60_398 VDD VSS sg13g2_decap_8
XFILLER_9_252 VDD VSS sg13g2_decap_8
Xclkload11 clkload11/Y _2365_/CLK VDD VSS sg13g2_inv_2
XFILLER_86_1055 VDD VSS sg13g2_decap_4
XFILLER_47_1006 VDD VSS sg13g2_decap_8
XFILLER_69_922 VDD VSS sg13g2_decap_8
X_1425_ _1424_/Y VDD _2233_/D VSS _1385_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_69_988 VDD VSS sg13g2_decap_8
XFILLER_29_819 VDD VSS sg13g2_decap_8
XFILLER_68_443 VDD VSS sg13g2_fill_1
X_1356_ _1357_/A _1347_/Y hold446/X _1347_/B _1379_/A VDD VSS sg13g2_a22oi_1
XFILLER_84_947 VDD VSS sg13g2_decap_8
XFILLER_96_796 VDD VSS sg13g2_decap_8
XFILLER_83_424 VDD VSS sg13g2_decap_8
XFILLER_23_1050 VDD VSS sg13g2_decap_8
XFILLER_56_616 VDD VSS sg13g2_decap_8
XFILLER_68_487 VDD VSS sg13g2_decap_8
XFILLER_28_329 VDD VSS sg13g2_decap_8
X_1287_ VDD _2173_/D _1287_/A VSS sg13g2_inv_1
XFILLER_49_690 VDD VSS sg13g2_decap_8
XFILLER_93_1004 VDD VSS sg13g2_decap_8
XFILLER_71_619 VDD VSS sg13g2_decap_8
XFILLER_37_896 VDD VSS sg13g2_decap_8
XFILLER_24_546 VDD VSS sg13g2_decap_8
XFILLER_34_28 VDD VSS sg13g2_decap_8
XFILLER_93_1059 VDD VSS sg13g2_fill_2
XFILLER_63_192 VDD VSS sg13g2_decap_8
Xclkload5 VDD clkload5/Y clkload5/A VSS sg13g2_inv_1
XFILLER_20_763 VDD VSS sg13g2_decap_8
XFILLER_30_1043 VDD VSS sg13g2_decap_8
XFILLER_3_406 VDD VSS sg13g2_decap_8
XFILLER_106_846 VDD VSS sg13g2_decap_8
XFILLER_79_708 VDD VSS sg13g2_decap_8
XFILLER_105_323 VDD VSS sg13g2_decap_8
XFILLER_59_14 VDD VSS sg13g2_decap_8
XFILLER_1_7 VDD VSS sg13g2_decap_8
XFILLER_99_590 VDD VSS sg13g2_decap_8
XFILLER_8_1022 VDD VSS sg13g2_decap_8
XFILLER_87_752 VDD VSS sg13g2_decap_8
XFILLER_59_465 VDD VSS sg13g2_fill_2
XFILLER_59_443 VDD VSS sg13g2_decap_4
XFILLER_75_936 VDD VSS sg13g2_decap_8
XFILLER_75_925 VDD VSS sg13g2_decap_8
XFILLER_101_573 VDD VSS sg13g2_decap_8
XFILLER_86_251 VDD VSS sg13g2_decap_8
XFILLER_74_424 VDD VSS sg13g2_decap_8
XFILLER_75_35 VDD VSS sg13g2_decap_8
XFILLER_47_616 VDD VSS sg13g2_decap_8
XFILLER_59_476 VDD VSS sg13g2_decap_8
XFILLER_19_329 VDD VSS sg13g2_decap_8
XFILLER_74_446 VDD VSS sg13g2_decap_8
XFILLER_74_468 VDD VSS sg13g2_decap_8
XFILLER_74_479 VDD VSS sg13g2_fill_2
XFILLER_43_800 VDD VSS sg13g2_decap_8
XFILLER_28_896 VDD VSS sg13g2_decap_8
XFILLER_91_56 VDD VSS sg13g2_decap_8
XFILLER_43_877 VDD VSS sg13g2_decap_8
XFILLER_15_546 VDD VSS sg13g2_decap_8
XFILLER_42_343 VDD VSS sg13g2_decap_8
XFILLER_70_696 VDD VSS sg13g2_decap_8
XFILLER_42_398 VDD VSS sg13g2_decap_8
XFILLER_11_763 VDD VSS sg13g2_decap_8
XFILLER_109_651 VDD VSS sg13g2_decap_8
XFILLER_10_273 VDD VSS sg13g2_decap_8
XFILLER_7_756 VDD VSS sg13g2_decap_8
XFILLER_108_161 VDD VSS sg13g2_decap_8
XFILLER_6_266 VDD VSS sg13g2_decap_8
XFILLER_112_805 VDD VSS sg13g2_decap_8
XFILLER_3_973 VDD VSS sg13g2_decap_8
XFILLER_97_549 VDD VSS sg13g2_decap_8
XFILLER_111_315 VDD VSS sg13g2_decap_8
XFILLER_69_218 VDD VSS sg13g2_decap_8
XFILLER_2_483 VDD VSS sg13g2_decap_8
XFILLER_34_7 VDD VSS sg13g2_decap_8
X_2190_ _2190_/RESET_B VSS VDD _2190_/D _2190_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_66_914 VDD VSS sg13g2_decap_8
X_1210_ VDD _1210_/Y _2249_/Q VSS sg13g2_inv_1
XFILLER_78_796 VDD VSS sg13g2_decap_4
XFILLER_77_273 VDD VSS sg13g2_decap_8
XFILLER_65_413 VDD VSS sg13g2_fill_2
XFILLER_1_21 VDD VSS sg13g2_decap_8
XFILLER_93_766 VDD VSS sg13g2_decap_8
XFILLER_92_221 VDD VSS sg13g2_decap_8
XFILLER_37_126 VDD VSS sg13g2_decap_8
XFILLER_81_939 VDD VSS sg13g2_decap_8
XFILLER_1_98 VDD VSS sg13g2_decap_8
XFILLER_92_298 VDD VSS sg13g2_decap_8
XFILLER_46_682 VDD VSS sg13g2_decap_8
XFILLER_34_833 VDD VSS sg13g2_decap_8
XFILLER_19_896 VDD VSS sg13g2_decap_8
XFILLER_60_140 VDD VSS sg13g2_decap_8
XFILLER_33_343 VDD VSS sg13g2_decap_8
X_1974_ _1973_/B _1973_/A _1973_/C _1974_/X VDD VSS sg13g2_a21o_1
XFILLER_53_1054 VDD VSS sg13g2_decap_8
XFILLER_60_0 VDD VSS sg13g2_decap_8
XFILLER_102_326 VDD VSS sg13g2_decap_8
XFILLER_69_741 VDD VSS sg13g2_decap_8
X_1408_ VDD _2226_/D _1408_/A VSS sg13g2_inv_1
XFILLER_29_28 VDD VSS sg13g2_decap_8
XFILLER_111_882 VDD VSS sg13g2_decap_8
XFILLER_96_571 VDD VSS sg13g2_decap_8
XFILLER_60_1025 VDD VSS sg13g2_decap_8
XFILLER_57_936 VDD VSS sg13g2_decap_8
XFILLER_29_616 VDD VSS sg13g2_decap_8
X_1339_ VDD _2199_/D _1339_/A VSS sg13g2_inv_1
XFILLER_84_733 VDD VSS sg13g2_decap_8
XFILLER_57_969 VDD VSS sg13g2_fill_1
XFILLER_68_284 VDD VSS sg13g2_decap_8
XFILLER_28_126 VDD VSS sg13g2_decap_8
XFILLER_84_788 VDD VSS sg13g2_decap_4
XFILLER_56_468 VDD VSS sg13g2_decap_4
XFILLER_37_693 VDD VSS sg13g2_decap_8
XFILLER_25_833 VDD VSS sg13g2_decap_8
XFILLER_45_49 VDD VSS sg13g2_decap_8
XFILLER_52_652 VDD VSS sg13g2_decap_4
XFILLER_24_343 VDD VSS sg13g2_decap_8
XFILLER_80_994 VDD VSS sg13g2_decap_8
XFILLER_51_140 VDD VSS sg13g2_fill_2
XFILLER_101_77 VDD VSS sg13g2_decap_8
XFILLER_40_858 VDD VSS sg13g2_decap_8
XFILLER_51_195 VDD VSS sg13g2_decap_8
XFILLER_20_560 VDD VSS sg13g2_decap_8
XFILLER_106_643 VDD VSS sg13g2_decap_8
XFILLER_3_203 VDD VSS sg13g2_decap_8
XFILLER_79_505 VDD VSS sg13g2_decap_8
XFILLER_10_63 VDD VSS sg13g2_decap_8
XFILLER_0_910 VDD VSS sg13g2_decap_8
X_2302__103 VDD VSS _2302_/RESET_B sg13g2_tiehi
XFILLER_86_56 VDD VSS sg13g2_decap_8
XFILLER_102_860 VDD VSS sg13g2_decap_8
XFILLER_75_700 VDD VSS sg13g2_decap_8
XFILLER_0_987 VDD VSS sg13g2_decap_8
XFILLER_59_284 VDD VSS sg13g2_decap_8
XFILLER_19_126 VDD VSS sg13g2_decap_8
XFILLER_47_435 VDD VSS sg13g2_decap_8
XFILLER_90_703 VDD VSS sg13g2_decap_8
XFILLER_74_265 VDD VSS sg13g2_decap_8
XFILLER_76_1010 VDD VSS sg13g2_fill_2
XFILLER_56_991 VDD VSS sg13g2_fill_1
XFILLER_28_693 VDD VSS sg13g2_decap_8
XFILLER_62_449 VDD VSS sg13g2_decap_8
XFILLER_16_833 VDD VSS sg13g2_decap_8
XFILLER_15_343 VDD VSS sg13g2_decap_8
XFILLER_43_674 VDD VSS sg13g2_decap_8
XFILLER_42_140 VDD VSS sg13g2_decap_8
XFILLER_42_151 VDD VSS sg13g2_fill_1
XFILLER_31_847 VDD VSS sg13g2_decap_8
XFILLER_42_184 VDD VSS sg13g2_decap_8
XFILLER_11_560 VDD VSS sg13g2_decap_8
XFILLER_30_357 VDD VSS sg13g2_decap_8
XFILLER_51_81 VDD VSS sg13g2_decap_8
X_1690_ _1725_/A _1690_/B _1690_/Y VDD VSS sg13g2_nor2_1
Xhold509 _1496_/Y VDD VSS _1497_/C sg13g2_dlygate4sd3_1
XFILLER_7_553 VDD VSS sg13g2_decap_8
XFILLER_100_1052 VDD VSS sg13g2_decap_8
XFILLER_112_602 VDD VSS sg13g2_decap_8
XFILLER_111_112 VDD VSS sg13g2_decap_8
X_2311_ _2311_/RESET_B VSS VDD _2311_/D _2311_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_3_770 VDD VSS sg13g2_decap_8
XFILLER_2_280 VDD VSS sg13g2_decap_8
XFILLER_112_679 VDD VSS sg13g2_decap_8
XFILLER_78_560 VDD VSS sg13g2_decap_4
X_2242_ _2242_/RESET_B VSS VDD _2242_/D _2242_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_97_379 VDD VSS sg13g2_decap_8
XFILLER_85_519 VDD VSS sg13g2_decap_8
XFILLER_66_722 VDD VSS sg13g2_decap_8
XFILLER_66_700 VDD VSS sg13g2_decap_8
X_2173_ _2173_/RESET_B VSS VDD _2173_/D _2173_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_111_189 VDD VSS sg13g2_decap_8
XFILLER_93_530 VDD VSS sg13g2_fill_2
XFILLER_39_969 VDD VSS sg13g2_decap_8
XFILLER_38_446 VDD VSS sg13g2_decap_8
XFILLER_93_563 VDD VSS sg13g2_decap_4
XFILLER_54_906 VDD VSS sg13g2_decap_8
XFILLER_65_254 VDD VSS sg13g2_fill_2
XFILLER_53_405 VDD VSS sg13g2_fill_1
XFILLER_81_736 VDD VSS sg13g2_decap_8
XFILLER_80_213 VDD VSS sg13g2_decap_8
XFILLER_65_276 VDD VSS sg13g2_fill_1
XFILLER_19_693 VDD VSS sg13g2_decap_8
XFILLER_34_630 VDD VSS sg13g2_decap_8
XFILLER_53_449 VDD VSS sg13g2_decap_8
XFILLER_90_1029 VDD VSS sg13g2_decap_8
XFILLER_61_460 VDD VSS sg13g2_decap_8
XFILLER_33_140 VDD VSS sg13g2_decap_8
XFILLER_22_847 VDD VSS sg13g2_decap_8
XFILLER_21_357 VDD VSS sg13g2_decap_8
X_1957_ VSS VDD _1982_/A _1958_/B _1958_/A sg13g2_or2_1
X_1888_ _1891_/A _1888_/A _1888_/B VDD VSS sg13g2_xnor2_1
XFILLER_1_707 VDD VSS sg13g2_decap_8
XFILLER_103_602 VDD VSS sg13g2_decap_8
XFILLER_0_217 VDD VSS sg13g2_decap_8
XFILLER_88_357 VDD VSS sg13g2_fill_2
XFILLER_88_346 VDD VSS sg13g2_decap_8
XFILLER_102_112 VDD VSS sg13g2_decap_8
XFILLER_103_679 VDD VSS sg13g2_decap_4
XFILLER_76_519 VDD VSS sg13g2_decap_8
XFILLER_69_593 VDD VSS sg13g2_decap_8
XFILLER_84_530 VDD VSS sg13g2_decap_8
XFILLER_57_744 VDD VSS sg13g2_decap_8
XFILLER_5_1036 VDD VSS sg13g2_decap_8
XFILLER_56_37 VDD VSS sg13g2_decap_8
XFILLER_29_413 VDD VSS sg13g2_decap_8
XFILLER_84_574 VDD VSS sg13g2_fill_2
XFILLER_84_563 VDD VSS sg13g2_decap_8
XFILLER_84_585 VDD VSS sg13g2_decap_8
XFILLER_112_21 VDD VSS sg13g2_decap_8
XFILLER_56_298 VDD VSS sg13g2_decap_8
XFILLER_72_14 VDD VSS sg13g2_decap_8
XFILLER_25_630 VDD VSS sg13g2_decap_8
XFILLER_37_490 VDD VSS sg13g2_decap_8
XFILLER_112_98 VDD VSS sg13g2_decap_8
XFILLER_53_983 VDD VSS sg13g2_decap_8
XFILLER_24_140 VDD VSS sg13g2_decap_8
XFILLER_13_847 VDD VSS sg13g2_decap_8
Xin_data_pads\[6\].in_data_pad IOVDD IOVSS _1385_/A in_data_PADs[6] VDD VSS sg13g2_IOPadIn
XFILLER_40_655 VDD VSS sg13g2_decap_8
XFILLER_12_357 VDD VSS sg13g2_decap_8
X_2189__162 VDD VSS _2189_/RESET_B sg13g2_tiehi
XFILLER_108_0 VDD VSS sg13g2_decap_8
XFILLER_4_567 VDD VSS sg13g2_decap_8
XFILLER_21_84 VDD VSS sg13g2_decap_8
XFILLER_107_996 VDD VSS sg13g2_decap_8
XFILLER_106_484 VDD VSS sg13g2_decap_4
XFILLER_79_313 VDD VSS sg13g2_decap_8
XFILLER_97_77 VDD VSS sg13g2_decap_8
XFILLER_43_1031 VDD VSS sg13g2_decap_8
XFILLER_0_784 VDD VSS sg13g2_decap_8
XFILLER_75_574 VDD VSS sg13g2_decap_8
XFILLER_36_917 VDD VSS sg13g2_decap_8
XFILLER_90_522 VDD VSS sg13g2_fill_2
XFILLER_90_511 VDD VSS sg13g2_decap_8
XFILLER_29_980 VDD VSS sg13g2_decap_8
XFILLER_46_70 VDD VSS sg13g2_decap_8
XFILLER_35_427 VDD VSS sg13g2_decap_8
XFILLER_63_758 VDD VSS sg13g2_decap_8
XFILLER_16_630 VDD VSS sg13g2_decap_8
XFILLER_28_490 VDD VSS sg13g2_decap_8
XFILLER_90_577 VDD VSS sg13g2_decap_4
XFILLER_15_140 VDD VSS sg13g2_decap_8
XFILLER_71_791 VDD VSS sg13g2_decap_8
XFILLER_31_644 VDD VSS sg13g2_decap_8
X_1811_ _1811_/B _1811_/A _1889_/A VDD VSS sg13g2_xor2_1
XFILLER_50_1002 VDD VSS sg13g2_decap_8
XFILLER_30_154 VDD VSS sg13g2_decap_8
XFILLER_62_91 VDD VSS sg13g2_decap_8
XFILLER_50_1024 VDD VSS sg13g2_decap_4
XFILLER_8_840 VDD VSS sg13g2_decap_8
X_1742_ _2241_/Q _2233_/Q _1772_/A VDD VSS sg13g2_xor2_1
XFILLER_7_350 VDD VSS sg13g2_decap_8
XFILLER_7_42 VDD VSS sg13g2_decap_8
XFILLER_11_1008 VDD VSS sg13g2_decap_8
Xhold306 _2190_/Q VDD VSS hold306/X sg13g2_dlygate4sd3_1
Xhold317 _1342_/Y VDD VSS _1343_/A sg13g2_dlygate4sd3_1
X_1673_ _1674_/A _1674_/B _1675_/B VDD VSS sg13g2_nor2_1
Xhold328 _1312_/Y VDD VSS _1313_/A sg13g2_dlygate4sd3_1
Xhold339 _1314_/Y VDD VSS _1315_/A sg13g2_dlygate4sd3_1
XFILLER_98_633 VDD VSS sg13g2_decap_8
Xout_data_pads\[7\].out_data_pad _2373_/Q IOVDD IOVSS out_data_PADs[7] VDD VSS sg13g2_IOPadOut30mA
XFILLER_100_616 VDD VSS sg13g2_decap_8
XFILLER_98_677 VDD VSS sg13g2_decap_8
XFILLER_112_476 VDD VSS sg13g2_decap_8
XFILLER_97_165 VDD VSS sg13g2_decap_8
XFILLER_23_0 VDD VSS sg13g2_decap_8
XFILLER_85_327 VDD VSS sg13g2_decap_8
X_2225_ _2225__90/L_HI VSS VDD _2225_/D _2225_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_38_210 VDD VSS sg13g2_decap_8
XFILLER_94_861 VDD VSS sg13g2_fill_1
XFILLER_27_917 VDD VSS sg13g2_decap_8
XFILLER_39_766 VDD VSS sg13g2_decap_8
X_2156_ _2156_/A _2040_/A _2335_/D VDD VSS sg13g2_nor2b_1
XFILLER_66_585 VDD VSS sg13g2_decap_8
XFILLER_26_427 VDD VSS sg13g2_decap_8
XFILLER_38_287 VDD VSS sg13g2_decap_8
XFILLER_81_566 VDD VSS sg13g2_fill_2
X_2087_ _2087_/Y _2065_/C _2089_/S _2062_/B _2004_/Y VDD VSS sg13g2_a22oi_1
XFILLER_54_758 VDD VSS sg13g2_decap_8
XFILLER_19_490 VDD VSS sg13g2_decap_8
X_2255__241 VDD VSS _2255_/RESET_B sg13g2_tiehi
Xclkbuf_leaf_18_clk clkbuf_leaf_0_clk/A _2289_/CLK VDD VSS sg13g2_buf_8
XFILLER_35_994 VDD VSS sg13g2_decap_8
XFILLER_107_1003 VDD VSS sg13g2_decap_8
XFILLER_50_953 VDD VSS sg13g2_decap_8
XFILLER_22_644 VDD VSS sg13g2_decap_8
XFILLER_21_154 VDD VSS sg13g2_decap_8
XFILLER_42_28 VDD VSS sg13g2_decap_8
XFILLER_108_738 VDD VSS sg13g2_decap_8
XFILLER_107_226 VDD VSS sg13g2_fill_2
XFILLER_107_215 VDD VSS sg13g2_fill_1
XFILLER_107_259 VDD VSS sg13g2_decap_8
XFILLER_101_7 VDD VSS sg13g2_decap_8
XFILLER_104_922 VDD VSS sg13g2_decap_8
XFILLER_107_21 VDD VSS sg13g2_decap_8
XFILLER_66_1042 VDD VSS sg13g2_decap_8
XFILLER_1_504 VDD VSS sg13g2_decap_8
XIO_CORNER_SOUTH_EAST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_103_421 VDD VSS sg13g2_fill_1
XFILLER_27_1015 VDD VSS sg13g2_decap_8
XFILLER_67_14 VDD VSS sg13g2_decap_8
XFILLER_104_999 VDD VSS sg13g2_decap_8
XFILLER_89_699 VDD VSS sg13g2_decap_8
XFILLER_103_465 VDD VSS sg13g2_fill_1
XFILLER_107_98 VDD VSS sg13g2_decap_8
XFILLER_88_154 VDD VSS sg13g2_decap_8
XFILLER_76_338 VDD VSS sg13g2_fill_2
XFILLER_29_210 VDD VSS sg13g2_decap_8
XFILLER_18_917 VDD VSS sg13g2_decap_8
XFILLER_72_522 VDD VSS sg13g2_decap_8
XFILLER_83_35 VDD VSS sg13g2_decap_8
XFILLER_57_574 VDD VSS sg13g2_decap_8
XFILLER_17_427 VDD VSS sg13g2_decap_8
XFILLER_29_287 VDD VSS sg13g2_decap_8
XFILLER_45_758 VDD VSS sg13g2_decap_8
XFILLER_72_577 VDD VSS sg13g2_decap_8
XFILLER_26_994 VDD VSS sg13g2_decap_8
XFILLER_44_257 VDD VSS sg13g2_decap_4
XFILLER_44_279 VDD VSS sg13g2_fill_1
XFILLER_16_84 VDD VSS sg13g2_decap_8
XFILLER_13_644 VDD VSS sg13g2_decap_8
XFILLER_41_986 VDD VSS sg13g2_decap_8
XFILLER_34_1008 VDD VSS sg13g2_decap_8
XFILLER_12_154 VDD VSS sg13g2_decap_8
XFILLER_9_637 VDD VSS sg13g2_decap_8
XFILLER_8_147 VDD VSS sg13g2_decap_8
XFILLER_5_854 VDD VSS sg13g2_decap_8
XFILLER_107_793 VDD VSS sg13g2_decap_8
XFILLER_99_419 VDD VSS sg13g2_fill_1
XFILLER_4_364 VDD VSS sg13g2_decap_8
XFILLER_110_914 VDD VSS sg13g2_decap_8
XFILLER_95_603 VDD VSS sg13g2_decap_8
XFILLER_95_614 VDD VSS sg13g2_fill_2
XFILLER_79_154 VDD VSS sg13g2_decap_8
XFILLER_95_658 VDD VSS sg13g2_decap_8
XFILLER_79_176 VDD VSS sg13g2_decap_8
XFILLER_0_581 VDD VSS sg13g2_decap_8
X_2010_ _2008_/X _2009_/X _2022_/S _2031_/A VDD VSS sg13g2_mux2_1
XFILLER_76_872 VDD VSS sg13g2_decap_8
XFILLER_48_596 VDD VSS sg13g2_decap_8
XFILLER_36_714 VDD VSS sg13g2_decap_8
XFILLER_91_864 VDD VSS sg13g2_fill_2
XFILLER_35_224 VDD VSS sg13g2_decap_8
XFILLER_63_588 VDD VSS sg13g2_fill_1
XFILLER_63_566 VDD VSS sg13g2_decap_8
XFILLER_51_717 VDD VSS sg13g2_decap_4
XFILLER_32_931 VDD VSS sg13g2_decap_8
XFILLER_17_994 VDD VSS sg13g2_decap_8
XFILLER_50_216 VDD VSS sg13g2_decap_8
XFILLER_50_238 VDD VSS sg13g2_decap_8
XFILLER_31_441 VDD VSS sg13g2_decap_8
X_1725_ _1725_/A _1724_/X _1725_/Y VDD VSS sg13g2_nor2b_1
Xclkbuf_leaf_7_clk clkbuf_leaf_9_clk/A _2371_/CLK VDD VSS sg13g2_buf_8
X_1656_ _1674_/B _2331_/Q _2323_/Q _2346_/Q _2338_/Q _2311_/Q _1656_/X VDD VSS sg13g2_mux4_1
X_1587_ _1595_/A _1587_/B _1587_/Y VDD VSS sg13g2_nor2_1
XFILLER_99_986 VDD VSS sg13g2_decap_8
XFILLER_101_914 VDD VSS sg13g2_decap_8
XFILLER_59_817 VDD VSS sg13g2_decap_8
XFILLER_86_658 VDD VSS sg13g2_fill_2
XFILLER_112_273 VDD VSS sg13g2_decap_8
XFILLER_58_316 VDD VSS sg13g2_decap_8
XFILLER_85_157 VDD VSS sg13g2_decap_8
XFILLER_37_28 VDD VSS sg13g2_decap_8
XFILLER_82_820 VDD VSS sg13g2_decap_8
XFILLER_39_563 VDD VSS sg13g2_decap_8
XFILLER_27_714 VDD VSS sg13g2_decap_8
XFILLER_66_371 VDD VSS sg13g2_decap_8
X_2208_ _2208_/RESET_B VSS VDD _2208_/D _2208_/Q clkload1/A sg13g2_dfrbpq_1
X_2139_ _2139_/A _2139_/B _2371_/D VDD VSS sg13g2_nor2_1
XFILLER_96_1046 VDD VSS sg13g2_decap_8
XFILLER_26_224 VDD VSS sg13g2_decap_8
X_2372__240 VDD VSS _2372_/RESET_B sg13g2_tiehi
XFILLER_82_886 VDD VSS sg13g2_decap_8
XFILLER_54_577 VDD VSS sg13g2_fill_2
XFILLER_42_728 VDD VSS sg13g2_decap_8
XFILLER_23_931 VDD VSS sg13g2_decap_8
XFILLER_35_791 VDD VSS sg13g2_decap_8
XFILLER_41_216 VDD VSS sg13g2_fill_2
XFILLER_22_441 VDD VSS sg13g2_decap_8
XFILLER_10_658 VDD VSS sg13g2_decap_8
XFILLER_108_535 VDD VSS sg13g2_decap_8
XFILLER_1_301 VDD VSS sg13g2_decap_8
XFILLER_78_35 VDD VSS sg13g2_decap_8
XFILLER_77_614 VDD VSS sg13g2_decap_8
XFILLER_89_474 VDD VSS sg13g2_fill_1
XFILLER_2_868 VDD VSS sg13g2_decap_8
XFILLER_104_785 VDD VSS sg13g2_decap_8
XFILLER_77_625 VDD VSS sg13g2_fill_2
XFILLER_103_284 VDD VSS sg13g2_decap_8
XFILLER_1_378 VDD VSS sg13g2_decap_8
XFILLER_49_316 VDD VSS sg13g2_decap_8
XFILLER_40_1012 VDD VSS sg13g2_decap_8
XFILLER_100_980 VDD VSS sg13g2_fill_2
XFILLER_92_628 VDD VSS sg13g2_decap_8
XFILLER_76_168 VDD VSS sg13g2_decap_8
XFILLER_94_56 VDD VSS sg13g2_decap_8
XFILLER_91_105 VDD VSS sg13g2_fill_2
XFILLER_18_714 VDD VSS sg13g2_decap_8
XFILLER_45_511 VDD VSS sg13g2_decap_8
XFILLER_73_853 VDD VSS sg13g2_decap_8
XFILLER_17_224 VDD VSS sg13g2_decap_8
XFILLER_72_352 VDD VSS sg13g2_decap_8
XFILLER_33_728 VDD VSS sg13g2_decap_8
XFILLER_60_503 VDD VSS sg13g2_decap_8
XFILLER_26_791 VDD VSS sg13g2_decap_8
XFILLER_14_931 VDD VSS sg13g2_decap_8
XFILLER_32_238 VDD VSS sg13g2_decap_8
XFILLER_13_441 VDD VSS sg13g2_decap_8
XFILLER_41_783 VDD VSS sg13g2_decap_8
XFILLER_9_434 VDD VSS sg13g2_decap_8
XFILLER_64_7 VDD VSS sg13g2_decap_8
XFILLER_99_205 VDD VSS sg13g2_decap_4
X_1510_ _1510_/B _2271_/Q _1510_/A _1516_/B VDD VSS sg13g2_nand3_1
XFILLER_5_651 VDD VSS sg13g2_decap_8
XFILLER_107_590 VDD VSS sg13g2_decap_8
X_1441_ VDD _2240_/D _1441_/A VSS sg13g2_inv_1
XFILLER_99_249 VDD VSS sg13g2_decap_8
XFILLER_4_21 VDD VSS sg13g2_decap_8
XFILLER_4_161 VDD VSS sg13g2_decap_8
XFILLER_110_711 VDD VSS sg13g2_decap_8
X_1372_ _1371_/Y VDD _2212_/D VSS _1367_/B _1370_/Y sg13g2_o21ai_1
XFILLER_4_98 VDD VSS sg13g2_decap_8
XFILLER_96_978 VDD VSS sg13g2_decap_8
XFILLER_95_455 VDD VSS sg13g2_decap_8
XFILLER_67_146 VDD VSS sg13g2_decap_8
XFILLER_110_788 VDD VSS sg13g2_decap_8
XFILLER_82_105 VDD VSS sg13g2_decap_4
XFILLER_49_883 VDD VSS sg13g2_decap_8
XFILLER_55_308 VDD VSS sg13g2_decap_8
XFILLER_36_511 VDD VSS sg13g2_decap_8
XFILLER_82_149 VDD VSS sg13g2_decap_8
XFILLER_36_588 VDD VSS sg13g2_decap_8
XFILLER_24_728 VDD VSS sg13g2_decap_8
XFILLER_63_352 VDD VSS sg13g2_decap_8
XFILLER_1_1050 VDD VSS sg13g2_decap_8
XFILLER_91_683 VDD VSS sg13g2_decap_8
XFILLER_90_160 VDD VSS sg13g2_decap_8
XFILLER_17_791 VDD VSS sg13g2_decap_8
XFILLER_23_238 VDD VSS sg13g2_decap_8
XFILLER_90_0 VDD VSS sg13g2_decap_8
XFILLER_51_558 VDD VSS sg13g2_decap_8
XFILLER_104_1006 VDD VSS sg13g2_decap_8
XFILLER_17_1036 VDD VSS sg13g2_decap_8
XFILLER_20_945 VDD VSS sg13g2_decap_8
X_1708_ _1714_/A _2317_/Q _2303_/Q VDD VSS sg13g2_xnor2_1
XFILLER_105_505 VDD VSS sg13g2_decap_8
X_1639_ _1639_/A _1638_/X _1639_/Y VDD VSS sg13g2_nor2b_1
XFILLER_63_1034 VDD VSS sg13g2_fill_1
XFILLER_87_956 VDD VSS sg13g2_decap_8
XFILLER_87_934 VDD VSS sg13g2_decap_8
XFILLER_101_733 VDD VSS sg13g2_decap_8
XFILLER_99_794 VDD VSS sg13g2_decap_8
XFILLER_98_260 VDD VSS sg13g2_decap_8
XFILLER_86_433 VDD VSS sg13g2_decap_8
XFILLER_48_49 VDD VSS sg13g2_decap_8
XFILLER_87_967 VDD VSS sg13g2_fill_1
XFILLER_74_606 VDD VSS sg13g2_decap_4
XFILLER_24_1029 VDD VSS sg13g2_decap_8
XFILLER_59_658 VDD VSS sg13g2_fill_2
XFILLER_58_135 VDD VSS sg13g2_decap_8
XFILLER_100_254 VDD VSS sg13g2_decap_8
XFILLER_73_105 VDD VSS sg13g2_decap_8
XFILLER_27_511 VDD VSS sg13g2_decap_8
XFILLER_46_319 VDD VSS sg13g2_decap_8
XFILLER_104_77 VDD VSS sg13g2_decap_8
XFILLER_67_691 VDD VSS sg13g2_decap_8
XFILLER_55_853 VDD VSS sg13g2_decap_8
XFILLER_70_801 VDD VSS sg13g2_decap_8
XFILLER_54_341 VDD VSS sg13g2_decap_8
XFILLER_15_728 VDD VSS sg13g2_decap_8
XFILLER_81_171 VDD VSS sg13g2_decap_4
XFILLER_27_588 VDD VSS sg13g2_decap_8
XFILLER_14_238 VDD VSS sg13g2_decap_8
Xfanout20 _1338_/B1 _1322_/B1 VDD VSS sg13g2_buf_1
XFILLER_70_878 VDD VSS sg13g2_decap_8
XFILLER_81_193 VDD VSS sg13g2_decap_4
XFILLER_80_14 VDD VSS sg13g2_decap_8
Xfanout31 _1346_/Y _1347_/B VDD VSS sg13g2_buf_1
Xfanout53 _1589_/C _1580_/A1 VDD VSS sg13g2_buf_1
Xfanout64 _1583_/A _1576_/A VDD VSS sg13g2_buf_1
Xfanout42 _1190_/Y _1527_/B VDD VSS sg13g2_buf_1
Xfanout75 _2138_/B1 _2150_/A VDD VSS sg13g2_buf_1
XFILLER_11_945 VDD VSS sg13g2_decap_8
XFILLER_109_833 VDD VSS sg13g2_decap_8
XFILLER_10_455 VDD VSS sg13g2_decap_8
XFILLER_13_63 VDD VSS sg13g2_decap_8
XFILLER_7_938 VDD VSS sg13g2_decap_8
XFILLER_6_448 VDD VSS sg13g2_decap_8
XFILLER_108_354 VDD VSS sg13g2_fill_2
XFILLER_89_56 VDD VSS sg13g2_decap_8
XFILLER_2_665 VDD VSS sg13g2_decap_8
XFILLER_78_923 VDD VSS sg13g2_decap_8
XFILLER_1_175 VDD VSS sg13g2_decap_8
XFILLER_89_293 VDD VSS sg13g2_decap_8
XFILLER_93_937 VDD VSS sg13g2_decap_8
XFILLER_92_403 VDD VSS sg13g2_fill_2
XFILLER_18_511 VDD VSS sg13g2_decap_8
XFILLER_37_308 VDD VSS sg13g2_decap_8
XFILLER_49_168 VDD VSS sg13g2_decap_8
XFILLER_46_831 VDD VSS sg13g2_decap_8
XFILLER_79_1052 VDD VSS sg13g2_decap_8
XFILLER_80_609 VDD VSS sg13g2_decap_8
XFILLER_72_182 VDD VSS sg13g2_decap_8
XFILLER_18_588 VDD VSS sg13g2_decap_8
XFILLER_33_525 VDD VSS sg13g2_decap_8
X_1990_ VSS VDD _2000_/A _1989_/Y _1990_/Y _2071_/B sg13g2_a21oi_1
XFILLER_54_92 VDD VSS sg13g2_decap_8
XFILLER_60_366 VDD VSS sg13g2_decap_4
XFILLER_9_231 VDD VSS sg13g2_decap_8
XFILLER_103_1050 VDD VSS sg13g2_decap_8
Xclkload12 _2371_/CLK clkload12/X VDD VSS sg13g2_buf_8
XFILLER_70_91 VDD VSS sg13g2_decap_8
XFILLER_87_208 VDD VSS sg13g2_decap_8
X_1424_ _1424_/Y _1424_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_69_978 VDD VSS sg13g2_fill_2
XFILLER_96_742 VDD VSS sg13g2_fill_2
XFILLER_95_241 VDD VSS sg13g2_decap_8
X_1355_ VDD _2206_/D _1355_/A VSS sg13g2_inv_1
XFILLER_84_937 VDD VSS sg13g2_fill_1
XFILLER_110_585 VDD VSS sg13g2_decap_8
XFILLER_96_775 VDD VSS sg13g2_decap_8
XFILLER_83_403 VDD VSS sg13g2_decap_8
XFILLER_68_466 VDD VSS sg13g2_decap_8
XFILLER_55_116 VDD VSS sg13g2_decap_8
XFILLER_28_308 VDD VSS sg13g2_decap_8
X_1286_ _1286_/Y _1344_/B1 hold310/X _1344_/A2 _2337_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_1054 VDD VSS sg13g2_decap_8
XFILLER_37_875 VDD VSS sg13g2_decap_8
XFILLER_70_119 VDD VSS sg13g2_decap_8
XFILLER_64_683 VDD VSS sg13g2_decap_8
XFILLER_24_525 VDD VSS sg13g2_decap_8
XFILLER_36_385 VDD VSS sg13g2_decap_8
XFILLER_52_856 VDD VSS sg13g2_decap_8
XFILLER_51_333 VDD VSS sg13g2_decap_8
XFILLER_51_388 VDD VSS sg13g2_decap_8
XFILLER_20_742 VDD VSS sg13g2_decap_8
Xclkload6 clkload6/A clkload6/X VDD VSS sg13g2_buf_8
XFILLER_50_28 VDD VSS sg13g2_fill_2
XFILLER_30_1022 VDD VSS sg13g2_decap_8
XFILLER_106_825 VDD VSS sg13g2_decap_8
XFILLER_105_302 VDD VSS sg13g2_decap_8
XFILLER_87_731 VDD VSS sg13g2_decap_8
XFILLER_105_379 VDD VSS sg13g2_decap_8
XFILLER_59_411 VDD VSS sg13g2_fill_2
XFILLER_8_1001 VDD VSS sg13g2_decap_8
XFILLER_101_541 VDD VSS sg13g2_decap_8
XFILLER_75_904 VDD VSS sg13g2_decap_8
XFILLER_86_230 VDD VSS sg13g2_decap_8
XFILLER_59_433 VDD VSS sg13g2_decap_4
XFILLER_86_274 VDD VSS sg13g2_decap_8
XFILLER_75_14 VDD VSS sg13g2_decap_8
XFILLER_19_308 VDD VSS sg13g2_decap_8
XFILLER_46_138 VDD VSS sg13g2_decap_8
XFILLER_28_875 VDD VSS sg13g2_decap_8
XFILLER_61_108 VDD VSS sg13g2_decap_8
XFILLER_83_981 VDD VSS sg13g2_fill_1
XFILLER_15_525 VDD VSS sg13g2_decap_8
XFILLER_27_385 VDD VSS sg13g2_decap_8
XFILLER_91_35 VDD VSS sg13g2_decap_8
XFILLER_43_856 VDD VSS sg13g2_decap_8
XFILLER_54_182 VDD VSS sg13g2_decap_8
XFILLER_70_675 VDD VSS sg13g2_decap_8
XFILLER_42_377 VDD VSS sg13g2_decap_8
X_2235__283 VDD VSS _2235_/RESET_B sg13g2_tiehi
XFILLER_11_742 VDD VSS sg13g2_decap_8
XFILLER_24_84 VDD VSS sg13g2_decap_8
XFILLER_30_539 VDD VSS sg13g2_decap_8
XFILLER_10_252 VDD VSS sg13g2_decap_8
XFILLER_109_630 VDD VSS sg13g2_decap_8
XFILLER_7_735 VDD VSS sg13g2_decap_8
XFILLER_108_140 VDD VSS sg13g2_decap_8
XFILLER_6_245 VDD VSS sg13g2_decap_8
XFILLER_97_517 VDD VSS sg13g2_fill_1
XFILLER_97_506 VDD VSS sg13g2_decap_8
XFILLER_3_952 VDD VSS sg13g2_decap_8
XFILLER_2_462 VDD VSS sg13g2_decap_8
XFILLER_27_7 VDD VSS sg13g2_decap_8
XFILLER_49_70 VDD VSS sg13g2_decap_4
X_2199__142 VDD VSS _2199_/RESET_B sg13g2_tiehi
XFILLER_78_775 VDD VSS sg13g2_decap_8
XFILLER_37_105 VDD VSS sg13g2_decap_8
XFILLER_93_745 VDD VSS sg13g2_decap_8
XFILLER_38_639 VDD VSS sg13g2_decap_8
XFILLER_81_918 VDD VSS sg13g2_fill_1
XFILLER_81_907 VDD VSS sg13g2_decap_8
XFILLER_53_609 VDD VSS sg13g2_decap_8
XFILLER_1_77 VDD VSS sg13g2_decap_8
XFILLER_19_875 VDD VSS sg13g2_decap_8
XFILLER_92_277 VDD VSS sg13g2_decap_8
XFILLER_80_439 VDD VSS sg13g2_decap_8
XFILLER_34_812 VDD VSS sg13g2_decap_8
XFILLER_18_385 VDD VSS sg13g2_decap_8
XFILLER_45_160 VDD VSS sg13g2_decap_4
XFILLER_65_80 VDD VSS sg13g2_decap_8
XFILLER_73_491 VDD VSS sg13g2_decap_8
XFILLER_33_322 VDD VSS sg13g2_decap_8
XFILLER_45_182 VDD VSS sg13g2_decap_8
XFILLER_92_1060 VDD VSS sg13g2_fill_1
XFILLER_53_1011 VDD VSS sg13g2_decap_8
XFILLER_61_697 VDD VSS sg13g2_fill_1
XFILLER_34_889 VDD VSS sg13g2_decap_8
X_1973_ _1973_/B _1973_/C _1973_/A _1973_/Y VDD VSS sg13g2_nand3_1
XFILLER_21_539 VDD VSS sg13g2_decap_8
XFILLER_33_399 VDD VSS sg13g2_decap_8
XFILLER_53_0 VDD VSS sg13g2_decap_8
XFILLER_88_517 VDD VSS sg13g2_decap_4
XFILLER_69_720 VDD VSS sg13g2_decap_8
X_1407_ _1408_/A _1392_/Y hold525/X _1391_/Y _1388_/A VDD VSS sg13g2_a22oi_1
XFILLER_60_1004 VDD VSS sg13g2_decap_8
XFILLER_111_861 VDD VSS sg13g2_decap_8
XFILLER_96_550 VDD VSS sg13g2_decap_8
XFILLER_69_797 VDD VSS sg13g2_decap_8
XFILLER_57_915 VDD VSS sg13g2_decap_8
XFILLER_28_105 VDD VSS sg13g2_decap_8
X_1338_ _1338_/Y _1338_/B1 hold399/X _1338_/A2 _2332_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_382 VDD VSS sg13g2_decap_8
XFILLER_83_222 VDD VSS sg13g2_fill_1
XFILLER_56_447 VDD VSS sg13g2_decap_8
X_1269_ VDD _2164_/D _1269_/A VSS sg13g2_inv_1
XFILLER_45_28 VDD VSS sg13g2_decap_8
XFILLER_83_299 VDD VSS sg13g2_decap_8
XFILLER_71_439 VDD VSS sg13g2_decap_8
XFILLER_37_672 VDD VSS sg13g2_decap_8
XFILLER_25_812 VDD VSS sg13g2_decap_8
XFILLER_43_119 VDD VSS sg13g2_decap_8
XFILLER_52_631 VDD VSS sg13g2_decap_8
XFILLER_24_322 VDD VSS sg13g2_decap_8
XFILLER_36_182 VDD VSS sg13g2_decap_8
XFILLER_80_973 VDD VSS sg13g2_decap_8
XFILLER_101_56 VDD VSS sg13g2_decap_8
XFILLER_40_837 VDD VSS sg13g2_decap_8
XFILLER_25_889 VDD VSS sg13g2_decap_8
XFILLER_12_539 VDD VSS sg13g2_decap_8
XFILLER_61_49 VDD VSS sg13g2_decap_8
XFILLER_24_399 VDD VSS sg13g2_decap_8
XFILLER_51_174 VDD VSS sg13g2_decap_8
XFILLER_106_622 VDD VSS sg13g2_decap_8
XFILLER_4_749 VDD VSS sg13g2_decap_8
XFILLER_3_259 VDD VSS sg13g2_decap_8
XFILLER_10_42 VDD VSS sg13g2_decap_8
XFILLER_106_699 VDD VSS sg13g2_decap_8
XFILLER_105_187 VDD VSS sg13g2_fill_1
XFILLER_86_35 VDD VSS sg13g2_decap_8
XFILLER_0_966 VDD VSS sg13g2_decap_8
XFILLER_48_937 VDD VSS sg13g2_decap_8
XFILLER_48_915 VDD VSS sg13g2_decap_4
XFILLER_59_252 VDD VSS sg13g2_fill_1
XFILLER_19_105 VDD VSS sg13g2_decap_8
XFILLER_47_414 VDD VSS sg13g2_fill_1
XFILLER_87_583 VDD VSS sg13g2_decap_8
XFILLER_75_756 VDD VSS sg13g2_decap_8
XFILLER_101_393 VDD VSS sg13g2_decap_8
XFILLER_59_274 VDD VSS sg13g2_fill_1
XFILLER_75_789 VDD VSS sg13g2_decap_8
XFILLER_74_244 VDD VSS sg13g2_decap_8
XFILLER_35_609 VDD VSS sg13g2_decap_8
XFILLER_19_84 VDD VSS sg13g2_decap_8
XFILLER_28_672 VDD VSS sg13g2_decap_8
XFILLER_62_428 VDD VSS sg13g2_decap_8
XFILLER_55_480 VDD VSS sg13g2_decap_8
XFILLER_16_812 VDD VSS sg13g2_decap_8
XFILLER_34_119 VDD VSS sg13g2_decap_8
XFILLER_76_1044 VDD VSS sg13g2_decap_8
XFILLER_90_759 VDD VSS sg13g2_decap_8
XFILLER_43_653 VDD VSS sg13g2_decap_8
XFILLER_15_322 VDD VSS sg13g2_decap_8
XFILLER_27_182 VDD VSS sg13g2_decap_8
XFILLER_71_984 VDD VSS sg13g2_decap_8
XFILLER_31_826 VDD VSS sg13g2_decap_8
XFILLER_16_889 VDD VSS sg13g2_decap_8
XFILLER_42_163 VDD VSS sg13g2_decap_8
XFILLER_15_399 VDD VSS sg13g2_decap_8
XFILLER_30_336 VDD VSS sg13g2_decap_8
XFILLER_7_532 VDD VSS sg13g2_decap_8
XFILLER_51_60 VDD VSS sg13g2_decap_8
XFILLER_13_1050 VDD VSS sg13g2_decap_8
XFILLER_83_1059 VDD VSS sg13g2_fill_2
XFILLER_98_848 VDD VSS sg13g2_fill_1
X_2310_ _2310_/RESET_B VSS VDD _2310_/D _2310_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_112_658 VDD VSS sg13g2_decap_8
X_2241_ _2241_/RESET_B VSS VDD _2241_/D _2241_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_97_336 VDD VSS sg13g2_decap_8
XFILLER_111_168 VDD VSS sg13g2_decap_8
XFILLER_39_948 VDD VSS sg13g2_decap_8
X_2172_ _2172_/RESET_B VSS VDD _2172_/D _2172_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_38_425 VDD VSS sg13g2_decap_8
XFILLER_81_715 VDD VSS sg13g2_decap_8
XFILLER_26_609 VDD VSS sg13g2_decap_8
XFILLER_65_233 VDD VSS sg13g2_decap_8
XFILLER_93_586 VDD VSS sg13g2_decap_8
XFILLER_47_992 VDD VSS sg13g2_decap_8
XFILLER_19_672 VDD VSS sg13g2_decap_8
XFILLER_20_1043 VDD VSS sg13g2_decap_8
XFILLER_25_119 VDD VSS sg13g2_decap_8
XFILLER_18_182 VDD VSS sg13g2_decap_8
XFILLER_90_1008 VDD VSS sg13g2_decap_8
XFILLER_80_269 VDD VSS sg13g2_decap_8
XFILLER_34_686 VDD VSS sg13g2_decap_8
XFILLER_22_826 VDD VSS sg13g2_decap_8
XFILLER_21_336 VDD VSS sg13g2_decap_8
XFILLER_33_196 VDD VSS sg13g2_decap_8
X_1956_ VSS VDD _1924_/A _1924_/B _1958_/B _1918_/X sg13g2_a21oi_1
X_1887_ _1887_/B _1887_/A _1967_/A VDD VSS sg13g2_xor2_1
XFILLER_88_325 VDD VSS sg13g2_decap_8
XFILLER_103_658 VDD VSS sg13g2_decap_8
XFILLER_89_859 VDD VSS sg13g2_decap_8
XFILLER_97_881 VDD VSS sg13g2_decap_8
XFILLER_69_572 VDD VSS sg13g2_decap_8
XFILLER_102_168 VDD VSS sg13g2_decap_8
XFILLER_99_1000 VDD VSS sg13g2_decap_8
XFILLER_57_723 VDD VSS sg13g2_decap_8
XFILLER_5_1015 VDD VSS sg13g2_decap_8
XFILLER_17_609 VDD VSS sg13g2_decap_8
XFILLER_29_469 VDD VSS sg13g2_decap_8
XIO_CORNER_NORTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_72_726 VDD VSS sg13g2_fill_1
XFILLER_56_277 VDD VSS sg13g2_decap_8
XFILLER_16_119 VDD VSS sg13g2_decap_8
XFILLER_44_439 VDD VSS sg13g2_decap_8
XFILLER_112_77 VDD VSS sg13g2_decap_8
XFILLER_53_962 VDD VSS sg13g2_decap_8
XFILLER_71_269 VDD VSS sg13g2_decap_8
XFILLER_25_686 VDD VSS sg13g2_decap_8
XFILLER_13_826 VDD VSS sg13g2_decap_8
XFILLER_80_781 VDD VSS sg13g2_decap_8
XFILLER_40_634 VDD VSS sg13g2_decap_8
XFILLER_12_336 VDD VSS sg13g2_decap_8
XFILLER_24_196 VDD VSS sg13g2_decap_8
XFILLER_36_1050 VDD VSS sg13g2_decap_8
XFILLER_9_819 VDD VSS sg13g2_decap_8
XFILLER_8_329 VDD VSS sg13g2_decap_8
XFILLER_21_63 VDD VSS sg13g2_decap_8
XFILLER_107_975 VDD VSS sg13g2_decap_8
XFILLER_4_546 VDD VSS sg13g2_decap_8
XFILLER_106_463 VDD VSS sg13g2_decap_8
XFILLER_97_56 VDD VSS sg13g2_decap_8
XFILLER_95_829 VDD VSS sg13g2_decap_8
XFILLER_94_317 VDD VSS sg13g2_decap_4
XFILLER_43_1010 VDD VSS sg13g2_decap_8
XFILLER_48_701 VDD VSS sg13g2_decap_8
XFILLER_0_763 VDD VSS sg13g2_decap_8
XFILLER_75_542 VDD VSS sg13g2_decap_8
XFILLER_63_737 VDD VSS sg13g2_decap_8
XFILLER_35_406 VDD VSS sg13g2_decap_8
XFILLER_90_556 VDD VSS sg13g2_decap_8
XFILLER_62_236 VDD VSS sg13g2_fill_1
XFILLER_47_299 VDD VSS sg13g2_fill_2
XFILLER_71_770 VDD VSS sg13g2_decap_8
XFILLER_44_984 VDD VSS sg13g2_decap_8
XFILLER_16_686 VDD VSS sg13g2_decap_8
XFILLER_50_409 VDD VSS sg13g2_decap_8
XFILLER_94_7 VDD VSS sg13g2_decap_8
XFILLER_31_623 VDD VSS sg13g2_decap_8
XFILLER_15_196 VDD VSS sg13g2_decap_8
X_1810_ _1801_/A VDD _1811_/B VSS _1812_/A _1812_/B sg13g2_o21ai_1
XFILLER_30_133 VDD VSS sg13g2_decap_8
XFILLER_62_70 VDD VSS sg13g2_decap_8
XFILLER_7_21 VDD VSS sg13g2_decap_8
X_1741_ _1741_/Y _2241_/Q _2233_/Q VDD VSS sg13g2_nand2b_1
Xhold307 _1320_/Y VDD VSS _1321_/A sg13g2_dlygate4sd3_1
X_1672_ _1681_/A _1688_/B _1641_/B VDD VSS sg13g2_nand2b_1
XFILLER_8_896 VDD VSS sg13g2_decap_8
Xhold318 _2171_/Q VDD VSS hold318/X sg13g2_dlygate4sd3_1
Xhold329 _2353_/Q VDD VSS _2102_/A sg13g2_dlygate4sd3_1
XFILLER_7_98 VDD VSS sg13g2_decap_8
XFILLER_98_612 VDD VSS sg13g2_decap_8
XFILLER_97_133 VDD VSS sg13g2_decap_8
XFILLER_112_455 VDD VSS sg13g2_decap_8
XFILLER_85_306 VDD VSS sg13g2_decap_8
XFILLER_79_881 VDD VSS sg13g2_decap_8
X_2224_ _2224__92/L_HI VSS VDD _2224_/D _2224_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_39_745 VDD VSS sg13g2_decap_8
X_2155_ _2156_/A _2040_/A _2334_/D VDD VSS sg13g2_nor2b_1
X_2359__277 VDD VSS _2359_/RESET_B sg13g2_tiehi
XFILLER_16_0 VDD VSS sg13g2_decap_8
XIO_BOND_in_data_pads\[5\].in_data_pad in_data_PADs[5] bondpad_70x70
XFILLER_93_383 VDD VSS sg13g2_decap_8
XFILLER_66_575 VDD VSS sg13g2_fill_1
XFILLER_53_203 VDD VSS sg13g2_decap_8
XFILLER_26_406 VDD VSS sg13g2_decap_8
XFILLER_38_266 VDD VSS sg13g2_decap_8
XFILLER_81_545 VDD VSS sg13g2_decap_8
X_2086_ _2086_/Y _2086_/A _2149_/A VDD VSS sg13g2_nand2_1
XFILLER_38_299 VDD VSS sg13g2_decap_8
XFILLER_35_973 VDD VSS sg13g2_decap_8
XFILLER_41_409 VDD VSS sg13g2_decap_8
XFILLER_50_932 VDD VSS sg13g2_decap_8
XFILLER_22_623 VDD VSS sg13g2_decap_8
XFILLER_61_280 VDD VSS sg13g2_decap_8
XFILLER_34_483 VDD VSS sg13g2_decap_8
XFILLER_21_133 VDD VSS sg13g2_decap_8
XFILLER_107_1059 VDD VSS sg13g2_fill_2
X_2331__185 VDD VSS _2331_/RESET_B sg13g2_tiehi
XFILLER_108_717 VDD VSS sg13g2_decap_8
X_1939_ _1940_/A _1939_/B _1939_/Y VDD VSS sg13g2_nor2_1
XFILLER_107_238 VDD VSS sg13g2_decap_8
XFILLER_104_901 VDD VSS sg13g2_decap_8
XFILLER_89_601 VDD VSS sg13g2_fill_1
XFILLER_66_1021 VDD VSS sg13g2_decap_8
XFILLER_89_645 VDD VSS sg13g2_decap_8
XFILLER_88_133 VDD VSS sg13g2_decap_8
XFILLER_104_978 VDD VSS sg13g2_decap_8
XFILLER_89_678 VDD VSS sg13g2_decap_8
XFILLER_103_444 VDD VSS sg13g2_decap_8
XFILLER_107_77 VDD VSS sg13g2_decap_8
XFILLER_45_704 VDD VSS sg13g2_decap_4
XFILLER_85_873 VDD VSS sg13g2_decap_8
XFILLER_83_14 VDD VSS sg13g2_decap_8
XFILLER_57_597 VDD VSS sg13g2_decap_8
XFILLER_45_737 VDD VSS sg13g2_decap_8
XFILLER_17_406 VDD VSS sg13g2_decap_8
XFILLER_29_266 VDD VSS sg13g2_decap_8
XFILLER_44_214 VDD VSS sg13g2_decap_8
XFILLER_44_225 VDD VSS sg13g2_fill_2
XFILLER_26_973 VDD VSS sg13g2_decap_8
XFILLER_60_729 VDD VSS sg13g2_decap_8
XFILLER_16_63 VDD VSS sg13g2_decap_8
XFILLER_13_623 VDD VSS sg13g2_decap_8
XFILLER_25_483 VDD VSS sg13g2_decap_8
XFILLER_73_1058 VDD VSS sg13g2_fill_2
XFILLER_41_965 VDD VSS sg13g2_decap_8
XFILLER_12_133 VDD VSS sg13g2_decap_8
XFILLER_9_616 VDD VSS sg13g2_decap_8
XFILLER_8_126 VDD VSS sg13g2_decap_8
XFILLER_5_833 VDD VSS sg13g2_decap_8
XFILLER_32_84 VDD VSS sg13g2_decap_8
XFILLER_4_343 VDD VSS sg13g2_decap_8
XFILLER_107_772 VDD VSS sg13g2_decap_8
XFILLER_79_133 VDD VSS sg13g2_decap_8
XFILLER_95_637 VDD VSS sg13g2_decap_4
XFILLER_0_560 VDD VSS sg13g2_decap_8
XFILLER_76_851 VDD VSS sg13g2_decap_8
XFILLER_94_147 VDD VSS sg13g2_decap_8
XFILLER_48_575 VDD VSS sg13g2_decap_8
XFILLER_57_81 VDD VSS sg13g2_decap_8
XFILLER_35_203 VDD VSS sg13g2_decap_8
XFILLER_63_545 VDD VSS sg13g2_decap_8
XFILLER_32_910 VDD VSS sg13g2_decap_8
XFILLER_17_973 VDD VSS sg13g2_decap_8
XFILLER_90_386 VDD VSS sg13g2_decap_8
XFILLER_73_91 VDD VSS sg13g2_decap_8
XFILLER_44_781 VDD VSS sg13g2_decap_8
XFILLER_16_483 VDD VSS sg13g2_decap_8
XFILLER_31_420 VDD VSS sg13g2_decap_8
X_2229__82 VDD VSS _2229__82/L_HI sg13g2_tiehi
XFILLER_32_987 VDD VSS sg13g2_decap_8
XFILLER_89_1010 VDD VSS sg13g2_decap_8
XFILLER_31_497 VDD VSS sg13g2_decap_8
XFILLER_89_1043 VDD VSS sg13g2_decap_8
X_1724_ hold559/X _1723_/Y _1724_/S _1724_/X VDD VSS sg13g2_mux2_1
XFILLER_8_693 VDD VSS sg13g2_decap_8
XFILLER_99_921 VDD VSS sg13g2_fill_2
X_1655_ _1671_/C _1655_/B _2301_/D VDD VSS sg13g2_nor2_1
XFILLER_99_965 VDD VSS sg13g2_decap_8
X_1586_ _1587_/B _1589_/A _1589_/C VDD VSS sg13g2_xnor2_1
XFILLER_112_252 VDD VSS sg13g2_decap_8
XFILLER_86_637 VDD VSS sg13g2_fill_2
XFILLER_100_425 VDD VSS sg13g2_decap_8
XFILLER_98_497 VDD VSS sg13g2_decap_8
XFILLER_39_520 VDD VSS sg13g2_fill_2
XFILLER_85_136 VDD VSS sg13g2_fill_1
X_2207_ _2207_/RESET_B VSS VDD _2207_/D _2207_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_2_1029 VDD VSS sg13g2_decap_8
XFILLER_26_203 VDD VSS sg13g2_decap_8
X_2138_ _2138_/B1 VDD _2139_/B VSS _2142_/A1 hold538/X sg13g2_o21ai_1
XFILLER_94_692 VDD VSS sg13g2_decap_8
XFILLER_82_865 VDD VSS sg13g2_decap_8
X_2069_ _1880_/Y _2086_/A _2069_/S _2069_/X VDD VSS sg13g2_mux2_1
XFILLER_54_589 VDD VSS sg13g2_decap_4
XFILLER_42_707 VDD VSS sg13g2_decap_8
XFILLER_35_770 VDD VSS sg13g2_decap_8
XFILLER_23_910 VDD VSS sg13g2_decap_8
XFILLER_22_420 VDD VSS sg13g2_decap_8
XFILLER_34_280 VDD VSS sg13g2_decap_8
XFILLER_23_987 VDD VSS sg13g2_decap_8
XFILLER_50_784 VDD VSS sg13g2_decap_8
XFILLER_10_637 VDD VSS sg13g2_decap_8
XFILLER_22_497 VDD VSS sg13g2_decap_8
XFILLER_78_14 VDD VSS sg13g2_decap_8
XFILLER_2_847 VDD VSS sg13g2_decap_8
XFILLER_104_764 VDD VSS sg13g2_decap_8
XFILLER_1_357 VDD VSS sg13g2_decap_8
XFILLER_103_263 VDD VSS sg13g2_decap_8
XFILLER_94_35 VDD VSS sg13g2_decap_8
XFILLER_76_147 VDD VSS sg13g2_decap_8
XFILLER_58_862 VDD VSS sg13g2_decap_8
XFILLER_17_203 VDD VSS sg13g2_decap_8
XFILLER_73_832 VDD VSS sg13g2_decap_8
XFILLER_84_191 VDD VSS sg13g2_decap_8
XFILLER_72_331 VDD VSS sg13g2_decap_8
XFILLER_57_383 VDD VSS sg13g2_decap_8
XFILLER_73_887 VDD VSS sg13g2_decap_8
XFILLER_45_567 VDD VSS sg13g2_decap_8
XFILLER_33_707 VDD VSS sg13g2_decap_8
XFILLER_27_84 VDD VSS sg13g2_decap_8
XFILLER_26_770 VDD VSS sg13g2_decap_8
XFILLER_14_910 VDD VSS sg13g2_decap_8
XFILLER_32_217 VDD VSS sg13g2_decap_8
XFILLER_60_559 VDD VSS sg13g2_decap_8
XFILLER_13_420 VDD VSS sg13g2_decap_8
XFILLER_25_280 VDD VSS sg13g2_decap_8
XFILLER_41_762 VDD VSS sg13g2_decap_8
XFILLER_9_413 VDD VSS sg13g2_decap_8
XFILLER_14_987 VDD VSS sg13g2_decap_8
XFILLER_13_497 VDD VSS sg13g2_decap_8
Xvss_pads\[0\].vss_pad IOVDD IOVSS VDD VSS sg13g2_IOPadVss
XFILLER_5_630 VDD VSS sg13g2_decap_8
XFILLER_4_140 VDD VSS sg13g2_decap_8
XFILLER_57_7 VDD VSS sg13g2_decap_8
X_1440_ _1441_/A _1429_/Y hold426/X _1429_/B _1382_/A VDD VSS sg13g2_a22oi_1
XFILLER_99_228 VDD VSS sg13g2_decap_8
XFILLER_49_1060 VDD VSS sg13g2_fill_1
XFILLER_96_913 VDD VSS sg13g2_decap_8
X_1371_ _1371_/Y _1371_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_4_77 VDD VSS sg13g2_decap_8
XFILLER_68_615 VDD VSS sg13g2_decap_8
XFILLER_110_767 VDD VSS sg13g2_decap_8
XFILLER_95_434 VDD VSS sg13g2_decap_8
XFILLER_68_659 VDD VSS sg13g2_decap_8
XFILLER_48_350 VDD VSS sg13g2_decap_8
XFILLER_76_692 VDD VSS sg13g2_decap_8
XFILLER_63_331 VDD VSS sg13g2_decap_8
XFILLER_91_651 VDD VSS sg13g2_decap_8
XFILLER_91_662 VDD VSS sg13g2_fill_2
XFILLER_64_887 VDD VSS sg13g2_decap_8
XFILLER_36_567 VDD VSS sg13g2_decap_8
XFILLER_24_707 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_51_537 VDD VSS sg13g2_decap_8
XFILLER_17_770 VDD VSS sg13g2_decap_8
XFILLER_23_217 VDD VSS sg13g2_decap_8
XFILLER_16_280 VDD VSS sg13g2_decap_8
XFILLER_17_1015 VDD VSS sg13g2_decap_8
XFILLER_32_784 VDD VSS sg13g2_decap_8
XFILLER_20_924 VDD VSS sg13g2_decap_8
XFILLER_83_0 VDD VSS sg13g2_decap_8
XFILLER_31_294 VDD VSS sg13g2_decap_8
XFILLER_9_980 VDD VSS sg13g2_decap_8
XFILLER_8_490 VDD VSS sg13g2_decap_8
X_1707_ _1725_/A _1707_/B _1707_/Y VDD VSS sg13g2_nor2_1
X_1638_ _2297_/Q _1637_/Y _1638_/S _1638_/X VDD VSS sg13g2_mux2_1
XFILLER_99_773 VDD VSS sg13g2_decap_8
XFILLER_86_412 VDD VSS sg13g2_decap_8
XFILLER_24_1008 VDD VSS sg13g2_decap_8
XFILLER_59_637 VDD VSS sg13g2_decap_8
XFILLER_48_28 VDD VSS sg13g2_decap_8
XFILLER_58_114 VDD VSS sg13g2_decap_8
X_1569_ _1576_/A _1569_/B _2280_/D VDD VSS sg13g2_nor2_1
XFILLER_86_489 VDD VSS sg13g2_decap_8
XFILLER_67_670 VDD VSS sg13g2_decap_8
XFILLER_104_56 VDD VSS sg13g2_decap_8
XFILLER_55_832 VDD VSS sg13g2_decap_8
XFILLER_54_320 VDD VSS sg13g2_decap_8
XFILLER_39_394 VDD VSS sg13g2_decap_8
XFILLER_27_567 VDD VSS sg13g2_decap_8
XFILLER_15_707 VDD VSS sg13g2_decap_8
XFILLER_64_49 VDD VSS sg13g2_decap_8
XFILLER_82_695 VDD VSS sg13g2_decap_8
XFILLER_81_150 VDD VSS sg13g2_decap_8
XFILLER_54_397 VDD VSS sg13g2_decap_8
XFILLER_14_217 VDD VSS sg13g2_decap_8
Xfanout21 fanout22/X _1338_/B1 VDD VSS sg13g2_buf_1
Xfanout10 _2036_/S _2061_/S VDD VSS sg13g2_buf_1
XFILLER_70_857 VDD VSS sg13g2_decap_8
Xfanout43 _1189_/Y _1671_/B VDD VSS sg13g2_buf_1
XFILLER_23_784 VDD VSS sg13g2_decap_8
Xfanout65 _1429_/A _1583_/A VDD VSS sg13g2_buf_1
Xfanout32 _1388_/B _1465_/C VDD VSS sg13g2_buf_1
XFILLER_11_924 VDD VSS sg13g2_decap_8
Xfanout54 _1577_/S0 _1589_/C VDD VSS sg13g2_buf_1
Xfanout76 _2138_/B1 _2071_/A VDD VSS sg13g2_buf_1
XFILLER_50_581 VDD VSS sg13g2_decap_8
XFILLER_50_592 VDD VSS sg13g2_fill_1
XFILLER_10_434 VDD VSS sg13g2_decap_8
XFILLER_13_42 VDD VSS sg13g2_decap_8
XFILLER_7_917 VDD VSS sg13g2_decap_8
XFILLER_22_294 VDD VSS sg13g2_decap_8
XFILLER_109_812 VDD VSS sg13g2_decap_8
XFILLER_6_427 VDD VSS sg13g2_decap_8
XFILLER_108_333 VDD VSS sg13g2_decap_8
XFILLER_109_889 VDD VSS sg13g2_decap_8
XFILLER_89_35 VDD VSS sg13g2_decap_8
XFILLER_78_902 VDD VSS sg13g2_decap_8
Xhold490 _2313_/Q VDD VSS hold490/X sg13g2_dlygate4sd3_1
XFILLER_2_644 VDD VSS sg13g2_decap_8
XFILLER_89_272 VDD VSS sg13g2_decap_8
XFILLER_77_412 VDD VSS sg13g2_decap_8
XFILLER_1_154 VDD VSS sg13g2_decap_8
XFILLER_49_103 VDD VSS sg13g2_decap_8
XFILLER_78_979 VDD VSS sg13g2_decap_8
XFILLER_77_445 VDD VSS sg13g2_fill_1
XFILLER_49_147 VDD VSS sg13g2_decap_8
XFILLER_77_489 VDD VSS sg13g2_decap_4
XFILLER_46_810 VDD VSS sg13g2_decap_8
XFILLER_64_106 VDD VSS sg13g2_decap_8
XFILLER_92_448 VDD VSS sg13g2_decap_8
XFILLER_64_117 VDD VSS sg13g2_fill_1
XFILLER_46_887 VDD VSS sg13g2_decap_8
XFILLER_46_854 VDD VSS sg13g2_fill_2
XFILLER_18_567 VDD VSS sg13g2_decap_8
XFILLER_33_504 VDD VSS sg13g2_decap_8
XFILLER_72_161 VDD VSS sg13g2_decap_8
XFILLER_61_879 VDD VSS sg13g2_decap_8
XFILLER_60_345 VDD VSS sg13g2_decap_8
XFILLER_54_71 VDD VSS sg13g2_decap_8
XFILLER_14_784 VDD VSS sg13g2_decap_8
XFILLER_13_294 VDD VSS sg13g2_decap_8
XFILLER_9_210 VDD VSS sg13g2_decap_8
XFILLER_70_70 VDD VSS sg13g2_decap_8
Xclkload13 VDD clkload13/Y _2369_/CLK VSS sg13g2_inv_1
XFILLER_9_287 VDD VSS sg13g2_decap_8
XFILLER_6_994 VDD VSS sg13g2_decap_8
XFILLER_102_509 VDD VSS sg13g2_fill_1
X_1423_ _1422_/Y VDD _2232_/D VSS _1382_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_96_721 VDD VSS sg13g2_decap_8
XFILLER_69_957 VDD VSS sg13g2_decap_8
XFILLER_96_754 VDD VSS sg13g2_decap_8
X_1354_ _1355_/A _1347_/Y hold455/X _1347_/B _1376_/A VDD VSS sg13g2_a22oi_1
XFILLER_68_434 VDD VSS sg13g2_decap_8
XFILLER_110_564 VDD VSS sg13g2_decap_8
X_1285_ VDD _2172_/D _1285_/A VSS sg13g2_inv_1
XFILLER_95_286 VDD VSS sg13g2_decap_8
XFILLER_110_1033 VDD VSS sg13g2_decap_8
XFILLER_92_960 VDD VSS sg13g2_decap_8
XFILLER_83_459 VDD VSS sg13g2_decap_8
XFILLER_64_662 VDD VSS sg13g2_decap_8
XFILLER_37_854 VDD VSS sg13g2_decap_8
XFILLER_52_824 VDD VSS sg13g2_decap_8
XFILLER_51_312 VDD VSS sg13g2_decap_8
XFILLER_24_504 VDD VSS sg13g2_decap_8
XFILLER_36_364 VDD VSS sg13g2_decap_8
XFILLER_32_581 VDD VSS sg13g2_decap_8
XFILLER_20_721 VDD VSS sg13g2_decap_8
Xclkload7 clkload7/A clkload7/Y VDD VSS sg13g2_inv_4
XFILLER_109_119 VDD VSS sg13g2_decap_8
XFILLER_30_1001 VDD VSS sg13g2_decap_8
XFILLER_20_798 VDD VSS sg13g2_decap_8
XFILLER_106_804 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[6\].out_data_pad out_data_PADs[6] bondpad_70x70
XFILLER_105_358 VDD VSS sg13g2_decap_8
XFILLER_87_710 VDD VSS sg13g2_decap_8
XFILLER_101_520 VDD VSS sg13g2_decap_8
XFILLER_8_1057 VDD VSS sg13g2_decap_4
XFILLER_87_787 VDD VSS sg13g2_decap_8
XIO_BOND_out_ready_pad out_ready_PAD bondpad_70x70
XFILLER_75_949 VDD VSS sg13g2_decap_8
XFILLER_46_117 VDD VSS sg13g2_decap_8
XFILLER_83_960 VDD VSS sg13g2_decap_8
XFILLER_55_662 VDD VSS sg13g2_decap_8
XFILLER_28_854 VDD VSS sg13g2_decap_8
XFILLER_83_993 VDD VSS sg13g2_decap_8
XFILLER_91_14 VDD VSS sg13g2_decap_8
XFILLER_43_835 VDD VSS sg13g2_decap_8
XFILLER_15_504 VDD VSS sg13g2_decap_8
XFILLER_54_150 VDD VSS sg13g2_fill_1
XFILLER_27_364 VDD VSS sg13g2_decap_8
XFILLER_42_301 VDD VSS sg13g2_decap_8
XFILLER_42_312 VDD VSS sg13g2_fill_2
XFILLER_70_654 VDD VSS sg13g2_decap_8
XFILLER_82_492 VDD VSS sg13g2_decap_8
XFILLER_30_518 VDD VSS sg13g2_decap_8
XFILLER_51_890 VDD VSS sg13g2_decap_8
XFILLER_23_581 VDD VSS sg13g2_decap_8
XFILLER_11_721 VDD VSS sg13g2_decap_8
XFILLER_24_63 VDD VSS sg13g2_decap_8
XFILLER_10_231 VDD VSS sg13g2_decap_8
XFILLER_7_714 VDD VSS sg13g2_decap_8
XFILLER_6_224 VDD VSS sg13g2_decap_8
XFILLER_11_798 VDD VSS sg13g2_decap_8
XFILLER_109_686 VDD VSS sg13g2_decap_8
XFILLER_3_931 VDD VSS sg13g2_decap_8
XFILLER_40_84 VDD VSS sg13g2_decap_8
XFILLER_2_441 VDD VSS sg13g2_decap_8
XFILLER_46_1052 VDD VSS sg13g2_decap_8
XFILLER_93_724 VDD VSS sg13g2_decap_8
XFILLER_77_242 VDD VSS sg13g2_decap_8
XFILLER_38_618 VDD VSS sg13g2_decap_8
XFILLER_66_949 VDD VSS sg13g2_decap_8
XFILLER_1_56 VDD VSS sg13g2_decap_8
XFILLER_92_256 VDD VSS sg13g2_decap_8
XFILLER_65_459 VDD VSS sg13g2_decap_8
XFILLER_19_854 VDD VSS sg13g2_decap_8
XFILLER_80_418 VDD VSS sg13g2_decap_8
XFILLER_73_470 VDD VSS sg13g2_decap_8
XFILLER_18_364 VDD VSS sg13g2_decap_8
XFILLER_45_150 VDD VSS sg13g2_fill_1
XFILLER_33_301 VDD VSS sg13g2_decap_8
XFILLER_34_868 VDD VSS sg13g2_decap_8
XFILLER_60_120 VDD VSS sg13g2_fill_1
XFILLER_21_518 VDD VSS sg13g2_decap_8
XFILLER_33_378 VDD VSS sg13g2_decap_8
X_1972_ _1973_/C _1972_/A _1972_/B VDD VSS sg13g2_xnor2_1
XFILLER_60_186 VDD VSS sg13g2_decap_8
XFILLER_14_581 VDD VSS sg13g2_decap_8
XFILLER_81_91 VDD VSS sg13g2_decap_8
XFILLER_14_1029 VDD VSS sg13g2_decap_8
XFILLER_6_791 VDD VSS sg13g2_decap_8
XFILLER_46_0 VDD VSS sg13g2_decap_8
XFILLER_103_829 VDD VSS sg13g2_decap_8
XFILLER_111_840 VDD VSS sg13g2_decap_8
X_1406_ VDD _2225_/D _1406_/A VSS sg13g2_inv_1
X_1337_ VDD _2198_/D _1337_/A VSS sg13g2_inv_1
XFILLER_69_776 VDD VSS sg13g2_decap_8
XFILLER_68_253 VDD VSS sg13g2_decap_8
XFILLER_68_264 VDD VSS sg13g2_fill_1
XFILLER_110_361 VDD VSS sg13g2_decap_8
XFILLER_56_426 VDD VSS sg13g2_decap_8
X_1268_ _1268_/Y _1280_/B1 hold394/X _1280_/A2 _2314_/Q VDD VSS sg13g2_a22oi_1
XFILLER_37_651 VDD VSS sg13g2_decap_8
XFILLER_83_278 VDD VSS sg13g2_decap_8
XFILLER_71_418 VDD VSS sg13g2_decap_8
X_1199_ VDD _1199_/Y _1199_/A VSS sg13g2_inv_1
XFILLER_52_610 VDD VSS sg13g2_decap_8
XFILLER_36_161 VDD VSS sg13g2_decap_8
XFILLER_24_301 VDD VSS sg13g2_decap_8
XFILLER_80_952 VDD VSS sg13g2_decap_8
XFILLER_25_868 VDD VSS sg13g2_decap_8
XFILLER_101_35 VDD VSS sg13g2_decap_8
XFILLER_52_665 VDD VSS sg13g2_fill_2
XFILLER_40_816 VDD VSS sg13g2_decap_8
XFILLER_12_518 VDD VSS sg13g2_decap_8
XFILLER_51_164 VDD VSS sg13g2_fill_2
XFILLER_24_378 VDD VSS sg13g2_decap_8
XFILLER_52_698 VDD VSS sg13g2_decap_8
XFILLER_61_28 VDD VSS sg13g2_decap_8
XFILLER_106_601 VDD VSS sg13g2_decap_8
XFILLER_20_595 VDD VSS sg13g2_decap_8
XFILLER_69_1052 VDD VSS sg13g2_decap_8
XFILLER_10_21 VDD VSS sg13g2_decap_8
XFILLER_4_728 VDD VSS sg13g2_decap_8
XFILLER_105_133 VDD VSS sg13g2_decap_8
XFILLER_3_238 VDD VSS sg13g2_decap_8
XFILLER_106_678 VDD VSS sg13g2_decap_8
XFILLER_86_14 VDD VSS sg13g2_decap_8
XFILLER_10_98 VDD VSS sg13g2_decap_8
XFILLER_0_945 VDD VSS sg13g2_decap_8
XFILLER_87_562 VDD VSS sg13g2_decap_8
XFILLER_102_895 VDD VSS sg13g2_decap_8
XFILLER_75_735 VDD VSS sg13g2_decap_8
XFILLER_101_372 VDD VSS sg13g2_decap_8
XFILLER_74_223 VDD VSS sg13g2_decap_8
XFILLER_19_63 VDD VSS sg13g2_decap_8
XFILLER_75_768 VDD VSS sg13g2_decap_8
XFILLER_28_651 VDD VSS sg13g2_decap_8
XFILLER_76_1012 VDD VSS sg13g2_fill_1
XFILLER_90_738 VDD VSS sg13g2_decap_8
XFILLER_62_407 VDD VSS sg13g2_decap_8
XFILLER_15_301 VDD VSS sg13g2_decap_8
XFILLER_27_161 VDD VSS sg13g2_decap_8
XFILLER_76_1034 VDD VSS sg13g2_fill_1
XFILLER_71_963 VDD VSS sg13g2_decap_8
XFILLER_43_632 VDD VSS sg13g2_decap_8
XFILLER_16_868 VDD VSS sg13g2_decap_8
XFILLER_37_1029 VDD VSS sg13g2_decap_8
XFILLER_31_805 VDD VSS sg13g2_decap_8
XFILLER_15_378 VDD VSS sg13g2_decap_8
XFILLER_35_84 VDD VSS sg13g2_decap_8
XFILLER_70_484 VDD VSS sg13g2_decap_8
XFILLER_30_315 VDD VSS sg13g2_decap_8
X_2313__267 VDD VSS _2313_/RESET_B sg13g2_tiehi
XFILLER_7_511 VDD VSS sg13g2_decap_8
XFILLER_11_595 VDD VSS sg13g2_decap_8
XFILLER_109_483 VDD VSS sg13g2_decap_8
XFILLER_7_588 VDD VSS sg13g2_decap_8
XFILLER_83_1038 VDD VSS sg13g2_decap_8
XFILLER_98_827 VDD VSS sg13g2_decap_8
XFILLER_97_315 VDD VSS sg13g2_decap_8
XFILLER_112_637 VDD VSS sg13g2_decap_8
X_2240_ _2240_/RESET_B VSS VDD _2240_/D _2240_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_111_147 VDD VSS sg13g2_decap_8
XFILLER_39_927 VDD VSS sg13g2_decap_8
XFILLER_38_404 VDD VSS sg13g2_decap_8
X_2171_ _2171_/RESET_B VSS VDD _2171_/D _2171_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_65_212 VDD VSS sg13g2_decap_8
XFILLER_93_554 VDD VSS sg13g2_decap_4
XFILLER_76_91 VDD VSS sg13g2_decap_8
XFILLER_66_768 VDD VSS sg13g2_decap_8
XFILLER_65_256 VDD VSS sg13g2_fill_1
XFILLER_19_651 VDD VSS sg13g2_decap_8
XFILLER_20_1022 VDD VSS sg13g2_decap_8
XFILLER_47_971 VDD VSS sg13g2_decap_8
XFILLER_18_161 VDD VSS sg13g2_decap_8
XFILLER_80_248 VDD VSS sg13g2_decap_8
XFILLER_62_974 VDD VSS sg13g2_decap_4
XFILLER_34_665 VDD VSS sg13g2_decap_8
XFILLER_22_805 VDD VSS sg13g2_decap_8
XFILLER_21_315 VDD VSS sg13g2_decap_8
XFILLER_33_175 VDD VSS sg13g2_decap_8
X_1955_ _1958_/A _1955_/A _1955_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_882 VDD VSS sg13g2_decap_8
X_1886_ _1972_/A _1972_/B _1886_/Y VDD VSS sg13g2_nor2_1
XFILLER_107_409 VDD VSS sg13g2_decap_8
XFILLER_88_304 VDD VSS sg13g2_decap_4
XFILLER_103_637 VDD VSS sg13g2_decap_8
XFILLER_97_860 VDD VSS sg13g2_decap_8
XFILLER_69_551 VDD VSS sg13g2_decap_8
XFILLER_102_147 VDD VSS sg13g2_decap_8
XFILLER_57_702 VDD VSS sg13g2_decap_8
XFILLER_99_1023 VDD VSS sg13g2_fill_2
X_2369_ _2369_/RESET_B VSS VDD _2369_/D _2369_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_84_510 VDD VSS sg13g2_decap_8
XFILLER_56_201 VDD VSS sg13g2_decap_8
XFILLER_56_28 VDD VSS sg13g2_decap_4
XFILLER_99_1056 VDD VSS sg13g2_decap_4
XFILLER_96_392 VDD VSS sg13g2_decap_8
XFILLER_45_919 VDD VSS sg13g2_decap_8
XFILLER_57_779 VDD VSS sg13g2_decap_8
XFILLER_56_256 VDD VSS sg13g2_decap_8
XFILLER_29_448 VDD VSS sg13g2_decap_8
XFILLER_38_982 VDD VSS sg13g2_decap_8
XFILLER_112_56 VDD VSS sg13g2_decap_8
XFILLER_80_760 VDD VSS sg13g2_decap_8
XFILLER_72_49 VDD VSS sg13g2_decap_8
XFILLER_25_665 VDD VSS sg13g2_decap_8
XFILLER_13_805 VDD VSS sg13g2_decap_8
XFILLER_40_613 VDD VSS sg13g2_decap_8
XFILLER_52_495 VDD VSS sg13g2_decap_4
XFILLER_12_315 VDD VSS sg13g2_decap_8
XFILLER_24_175 VDD VSS sg13g2_decap_8
XFILLER_8_308 VDD VSS sg13g2_decap_8
XFILLER_21_882 VDD VSS sg13g2_decap_8
XFILLER_20_392 VDD VSS sg13g2_decap_8
XFILLER_4_525 VDD VSS sg13g2_decap_8
XFILLER_21_42 VDD VSS sg13g2_decap_8
XFILLER_107_954 VDD VSS sg13g2_decap_8
XFILLER_106_442 VDD VSS sg13g2_decap_8
XFILLER_97_35 VDD VSS sg13g2_decap_8
XFILLER_79_348 VDD VSS sg13g2_decap_8
XFILLER_95_808 VDD VSS sg13g2_decap_8
XFILLER_79_359 VDD VSS sg13g2_fill_1
XFILLER_0_742 VDD VSS sg13g2_decap_8
XFILLER_88_893 VDD VSS sg13g2_decap_8
XFILLER_87_381 VDD VSS sg13g2_decap_8
XFILLER_75_521 VDD VSS sg13g2_decap_8
XFILLER_47_212 VDD VSS sg13g2_fill_1
XFILLER_48_768 VDD VSS sg13g2_decap_8
XFILLER_47_245 VDD VSS sg13g2_fill_1
XFILLER_63_716 VDD VSS sg13g2_decap_8
XFILLER_47_278 VDD VSS sg13g2_decap_8
XFILLER_90_535 VDD VSS sg13g2_decap_8
XFILLER_44_963 VDD VSS sg13g2_decap_8
XFILLER_31_602 VDD VSS sg13g2_decap_8
XFILLER_16_665 VDD VSS sg13g2_decap_8
XFILLER_43_462 VDD VSS sg13g2_decap_8
XFILLER_15_175 VDD VSS sg13g2_decap_8
XFILLER_30_112 VDD VSS sg13g2_decap_8
XFILLER_70_292 VDD VSS sg13g2_decap_8
XFILLER_87_7 VDD VSS sg13g2_decap_8
XFILLER_31_679 VDD VSS sg13g2_decap_8
XFILLER_12_882 VDD VSS sg13g2_decap_8
X_2168__204 VDD VSS _2168_/RESET_B sg13g2_tiehi
X_1740_ _2242_/Q _2234_/Q _1774_/A VDD VSS sg13g2_xor2_1
XFILLER_50_1059 VDD VSS sg13g2_fill_2
XFILLER_11_392 VDD VSS sg13g2_decap_8
XFILLER_30_189 VDD VSS sg13g2_decap_8
Xhold308 _2180_/Q VDD VSS hold308/X sg13g2_dlygate4sd3_1
X_1671_ _1680_/A _1671_/B _1671_/C _1671_/D _2309_/D VDD VSS sg13g2_nor4_1
XFILLER_7_77 VDD VSS sg13g2_decap_8
XFILLER_8_875 VDD VSS sg13g2_decap_8
Xhold319 _1282_/Y VDD VSS _1283_/A sg13g2_dlygate4sd3_1
XFILLER_7_385 VDD VSS sg13g2_decap_8
XFILLER_98_602 VDD VSS sg13g2_decap_4
XFILLER_112_434 VDD VSS sg13g2_decap_8
XFILLER_97_112 VDD VSS sg13g2_decap_8
XFILLER_97_156 VDD VSS sg13g2_fill_2
X_2223_ _2223__94/L_HI VSS VDD _2223_/D _2223_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_39_724 VDD VSS sg13g2_decap_8
X_2154_ _2162_/B _1826_/B _2333_/D VDD VSS sg13g2_nor2b_1
XFILLER_66_554 VDD VSS sg13g2_decap_8
XFILLER_38_245 VDD VSS sg13g2_decap_8
XFILLER_94_885 VDD VSS sg13g2_decap_8
XFILLER_93_362 VDD VSS sg13g2_decap_8
XFILLER_54_705 VDD VSS sg13g2_decap_8
XFILLER_81_524 VDD VSS sg13g2_decap_8
X_2085_ _2086_/A _2149_/A _2085_/X VDD VSS sg13g2_and2_1
XFILLER_81_568 VDD VSS sg13g2_fill_1
XFILLER_35_952 VDD VSS sg13g2_decap_8
XFILLER_50_911 VDD VSS sg13g2_decap_8
XFILLER_22_602 VDD VSS sg13g2_decap_8
XFILLER_62_782 VDD VSS sg13g2_decap_8
XFILLER_21_112 VDD VSS sg13g2_decap_8
XFILLER_34_462 VDD VSS sg13g2_decap_8
XFILLER_107_1038 VDD VSS sg13g2_decap_8
XFILLER_50_988 VDD VSS sg13g2_decap_8
XFILLER_22_679 VDD VSS sg13g2_decap_8
XFILLER_10_819 VDD VSS sg13g2_decap_8
X_1938_ _1938_/B _1938_/A _1992_/A VDD VSS sg13g2_xor2_1
XFILLER_21_189 VDD VSS sg13g2_decap_8
XFILLER_107_228 VDD VSS sg13g2_fill_1
X_1869_ _1869_/A _1869_/B _1870_/B VDD VSS sg13g2_and2_1
XFILLER_66_1000 VDD VSS sg13g2_decap_8
XFILLER_104_957 VDD VSS sg13g2_decap_8
XFILLER_89_624 VDD VSS sg13g2_decap_8
XFILLER_107_56 VDD VSS sg13g2_decap_8
XFILLER_88_112 VDD VSS sg13g2_decap_8
XFILLER_1_539 VDD VSS sg13g2_decap_8
XFILLER_103_489 VDD VSS sg13g2_decap_8
XFILLER_57_521 VDD VSS sg13g2_decap_8
XFILLER_67_49 VDD VSS sg13g2_decap_8
XFILLER_29_245 VDD VSS sg13g2_decap_8
XFILLER_84_362 VDD VSS sg13g2_decap_8
XFILLER_72_557 VDD VSS sg13g2_fill_2
XFILLER_26_952 VDD VSS sg13g2_decap_8
XFILLER_16_42 VDD VSS sg13g2_decap_8
XFILLER_44_248 VDD VSS sg13g2_decap_4
XFILLER_73_1037 VDD VSS sg13g2_decap_8
XFILLER_41_944 VDD VSS sg13g2_decap_8
XFILLER_13_602 VDD VSS sg13g2_decap_8
XFILLER_25_462 VDD VSS sg13g2_decap_8
XFILLER_12_112 VDD VSS sg13g2_decap_8
XFILLER_40_454 VDD VSS sg13g2_decap_8
XFILLER_52_281 VDD VSS sg13g2_fill_2
XFILLER_8_105 VDD VSS sg13g2_decap_8
XFILLER_13_679 VDD VSS sg13g2_decap_8
XFILLER_12_189 VDD VSS sg13g2_decap_8
XFILLER_32_63 VDD VSS sg13g2_decap_8
XFILLER_40_498 VDD VSS sg13g2_decap_8
XFILLER_5_812 VDD VSS sg13g2_decap_8
XFILLER_4_322 VDD VSS sg13g2_decap_8
XFILLER_10_1043 VDD VSS sg13g2_decap_8
XFILLER_107_751 VDD VSS sg13g2_decap_8
XFILLER_5_889 VDD VSS sg13g2_decap_8
XFILLER_79_112 VDD VSS sg13g2_decap_8
XFILLER_4_399 VDD VSS sg13g2_decap_8
XFILLER_80_1008 VDD VSS sg13g2_decap_8
XFILLER_110_949 VDD VSS sg13g2_decap_8
XFILLER_94_126 VDD VSS sg13g2_decap_8
XFILLER_67_329 VDD VSS sg13g2_decap_8
XFILLER_48_510 VDD VSS sg13g2_decap_8
XFILLER_76_830 VDD VSS sg13g2_decap_8
XFILLER_57_60 VDD VSS sg13g2_decap_8
XFILLER_91_822 VDD VSS sg13g2_decap_4
XFILLER_75_362 VDD VSS sg13g2_fill_1
XFILLER_36_749 VDD VSS sg13g2_decap_8
XFILLER_63_524 VDD VSS sg13g2_decap_8
XFILLER_91_866 VDD VSS sg13g2_fill_1
XFILLER_44_760 VDD VSS sg13g2_decap_8
XFILLER_17_952 VDD VSS sg13g2_decap_8
XFILLER_35_259 VDD VSS sg13g2_decap_8
XFILLER_73_70 VDD VSS sg13g2_decap_8
XFILLER_16_462 VDD VSS sg13g2_decap_8
XFILLER_32_966 VDD VSS sg13g2_decap_8
XFILLER_43_292 VDD VSS sg13g2_decap_8
XFILLER_43_281 VDD VSS sg13g2_fill_1
XFILLER_31_476 VDD VSS sg13g2_decap_8
XFILLER_106_1060 VDD VSS sg13g2_fill_1
X_1723_ _1723_/Y _1723_/A _1723_/B VDD VSS sg13g2_xnor2_1
XFILLER_8_672 VDD VSS sg13g2_decap_8
XFILLER_7_182 VDD VSS sg13g2_decap_8
X_1654_ _1654_/Y _1646_/Y _1653_/X _1697_/B _1671_/B VDD VSS sg13g2_a22oi_1
XFILLER_99_911 VDD VSS sg13g2_fill_1
XFILLER_104_209 VDD VSS sg13g2_decap_4
XFILLER_98_432 VDD VSS sg13g2_decap_8
X_1585_ _1595_/A _1602_/B _1521_/B VDD VSS sg13g2_nand2b_1
XFILLER_112_231 VDD VSS sg13g2_decap_8
XFILLER_101_949 VDD VSS sg13g2_decap_8
XFILLER_86_649 VDD VSS sg13g2_fill_2
XFILLER_98_476 VDD VSS sg13g2_decap_8
XFILLER_85_115 VDD VSS sg13g2_decap_8
XFILLER_26_1050 VDD VSS sg13g2_decap_8
XFILLER_100_448 VDD VSS sg13g2_decap_8
X_2206_ _2206_/RESET_B VSS VDD _2206_/D _2206_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_67_841 VDD VSS sg13g2_decap_8
XFILLER_67_896 VDD VSS sg13g2_decap_8
XFILLER_66_362 VDD VSS sg13g2_decap_4
XFILLER_66_340 VDD VSS sg13g2_fill_2
XFILLER_54_502 VDD VSS sg13g2_decap_8
XFILLER_2_1008 VDD VSS sg13g2_decap_8
X_2137_ VDD VSS _1206_/Y _2120_/A _2136_/X hold302/X _2139_/A _2124_/Y sg13g2_a221oi_1
XFILLER_82_855 VDD VSS sg13g2_decap_4
XFILLER_39_598 VDD VSS sg13g2_decap_8
XFILLER_27_749 VDD VSS sg13g2_decap_8
X_2068_ _2072_/A _2068_/B _2025_/A VDD VSS sg13g2_nand2b_1
XFILLER_53_18 VDD VSS sg13g2_fill_1
XFILLER_26_259 VDD VSS sg13g2_decap_8
XFILLER_81_398 VDD VSS sg13g2_decap_8
XFILLER_41_218 VDD VSS sg13g2_fill_1
Xout_data_pads\[3\].out_data_pad _2369_/Q IOVDD IOVSS out_data_PADs[3] VDD VSS sg13g2_IOPadOut30mA
XFILLER_23_966 VDD VSS sg13g2_decap_8
XFILLER_50_763 VDD VSS sg13g2_decap_8
XFILLER_10_616 VDD VSS sg13g2_decap_8
XFILLER_22_476 VDD VSS sg13g2_decap_8
XFILLER_33_1043 VDD VSS sg13g2_decap_8
XFILLER_6_609 VDD VSS sg13g2_decap_8
XFILLER_108_515 VDD VSS sg13g2_fill_1
XFILLER_5_119 VDD VSS sg13g2_decap_8
XFILLER_104_710 VDD VSS sg13g2_decap_8
XFILLER_2_826 VDD VSS sg13g2_decap_8
XFILLER_104_743 VDD VSS sg13g2_decap_8
XFILLER_103_242 VDD VSS sg13g2_decap_8
XFILLER_1_336 VDD VSS sg13g2_decap_8
XFILLER_89_487 VDD VSS sg13g2_decap_8
XFILLER_94_14 VDD VSS sg13g2_decap_8
XFILLER_76_126 VDD VSS sg13g2_decap_8
XFILLER_58_830 VDD VSS sg13g2_fill_1
XFILLER_100_982 VDD VSS sg13g2_fill_1
XFILLER_91_107 VDD VSS sg13g2_fill_1
XFILLER_40_1047 VDD VSS sg13g2_decap_8
XFILLER_85_682 VDD VSS sg13g2_decap_8
XFILLER_84_170 VDD VSS sg13g2_decap_8
XFILLER_45_546 VDD VSS sg13g2_decap_8
XFILLER_18_749 VDD VSS sg13g2_decap_8
XFILLER_27_63 VDD VSS sg13g2_decap_8
XFILLER_17_259 VDD VSS sg13g2_decap_8
XFILLER_72_387 VDD VSS sg13g2_decap_4
XFILLER_60_538 VDD VSS sg13g2_decap_8
XFILLER_41_741 VDD VSS sg13g2_decap_8
XFILLER_14_966 VDD VSS sg13g2_decap_8
XFILLER_13_476 VDD VSS sg13g2_decap_8
XFILLER_43_84 VDD VSS sg13g2_decap_8
XFILLER_9_469 VDD VSS sg13g2_decap_8
XFILLER_5_686 VDD VSS sg13g2_decap_8
X_1370_ _1370_/Y _1370_/A _1465_/C VDD VSS sg13g2_nand2_1
XFILLER_4_196 VDD VSS sg13g2_decap_8
XFILLER_4_56 VDD VSS sg13g2_decap_8
XFILLER_96_947 VDD VSS sg13g2_decap_8
XFILLER_95_413 VDD VSS sg13g2_decap_8
XFILLER_110_746 VDD VSS sg13g2_decap_8
XFILLER_67_126 VDD VSS sg13g2_fill_2
XFILLER_83_619 VDD VSS sg13g2_decap_8
XFILLER_76_671 VDD VSS sg13g2_decap_8
XFILLER_49_863 VDD VSS sg13g2_decap_4
XFILLER_91_630 VDD VSS sg13g2_decap_8
XFILLER_64_844 VDD VSS sg13g2_decap_8
XFILLER_48_395 VDD VSS sg13g2_decap_8
XFILLER_75_192 VDD VSS sg13g2_decap_8
XFILLER_84_91 VDD VSS sg13g2_decap_8
XFILLER_64_866 VDD VSS sg13g2_decap_8
XFILLER_36_546 VDD VSS sg13g2_decap_8
XFILLER_56_1010 VDD VSS sg13g2_fill_2
XFILLER_63_387 VDD VSS sg13g2_decap_8
XFILLER_90_195 VDD VSS sg13g2_decap_8
XFILLER_56_1043 VDD VSS sg13g2_decap_8
XFILLER_32_763 VDD VSS sg13g2_decap_8
XFILLER_20_903 VDD VSS sg13g2_decap_8
XFILLER_31_273 VDD VSS sg13g2_decap_8
XFILLER_76_0 VDD VSS sg13g2_decap_8
X_1706_ _1705_/Y VDD _1707_/B VSS _1720_/A hold506/X sg13g2_o21ai_1
X_1637_ _1637_/Y _1637_/A _1637_/B VDD VSS sg13g2_xnor2_1
XFILLER_87_903 VDD VSS sg13g2_decap_8
XFILLER_63_1014 VDD VSS sg13g2_fill_1
XFILLER_63_1003 VDD VSS sg13g2_decap_8
XFILLER_101_713 VDD VSS sg13g2_decap_8
XFILLER_63_1058 VDD VSS sg13g2_fill_2
XFILLER_59_616 VDD VSS sg13g2_decap_8
X_1568_ _1568_/Y _1527_/Y _1567_/Y hold463/X _1527_/B VDD VSS sg13g2_a22oi_1
X_1499_ VSS VDD hold295/X _1497_/B _1499_/Y _1498_/Y sg13g2_a21oi_1
XFILLER_95_980 VDD VSS sg13g2_decap_8
XFILLER_101_779 VDD VSS sg13g2_decap_8
XFILLER_86_468 VDD VSS sg13g2_decap_8
XFILLER_104_35 VDD VSS sg13g2_decap_8
XFILLER_55_811 VDD VSS sg13g2_decap_8
XFILLER_66_181 VDD VSS sg13g2_decap_8
XFILLER_39_373 VDD VSS sg13g2_decap_8
XFILLER_27_546 VDD VSS sg13g2_decap_8
XFILLER_64_28 VDD VSS sg13g2_decap_8
XFILLER_82_674 VDD VSS sg13g2_decap_8
XFILLER_70_836 VDD VSS sg13g2_decap_8
XFILLER_55_888 VDD VSS sg13g2_decap_8
Xfanout11 _2036_/S _2022_/S VDD VSS sg13g2_buf_1
Xfanout22 _1265_/X fanout22/X VDD VSS sg13g2_buf_1
XFILLER_70_1018 VDD VSS sg13g2_fill_2
Xfanout55 _1577_/S0 _1556_/S0 VDD VSS sg13g2_buf_1
Xfanout44 _2356_/Q _1259_/A VDD VSS sg13g2_buf_1
XFILLER_50_560 VDD VSS sg13g2_decap_8
XFILLER_23_763 VDD VSS sg13g2_decap_8
XFILLER_11_903 VDD VSS sg13g2_decap_8
Xfanout33 _1522_/Y _1523_/B VDD VSS sg13g2_buf_1
XFILLER_70_1029 VDD VSS sg13g2_fill_1
XFILLER_80_49 VDD VSS sg13g2_decap_8
Xfanout77 _2138_/B1 _1688_/B VDD VSS sg13g2_buf_1
Xfanout66 _2101_/A _1429_/A VDD VSS sg13g2_buf_1
XFILLER_10_413 VDD VSS sg13g2_decap_8
XFILLER_13_21 VDD VSS sg13g2_decap_8
XFILLER_22_273 VDD VSS sg13g2_decap_8
XFILLER_6_406 VDD VSS sg13g2_decap_8
XFILLER_108_312 VDD VSS sg13g2_fill_2
XFILLER_89_14 VDD VSS sg13g2_decap_8
XFILLER_13_98 VDD VSS sg13g2_decap_8
XFILLER_109_868 VDD VSS sg13g2_decap_8
XFILLER_108_356 VDD VSS sg13g2_fill_1
XFILLER_2_623 VDD VSS sg13g2_decap_8
Xhold480 _2241_/Q VDD VSS hold480/X sg13g2_dlygate4sd3_1
XFILLER_1_133 VDD VSS sg13g2_decap_8
XFILLER_104_584 VDD VSS sg13g2_decap_8
XFILLER_89_251 VDD VSS sg13g2_decap_8
Xhold491 _1689_/Y VDD VSS _1690_/B sg13g2_dlygate4sd3_1
XFILLER_78_958 VDD VSS sg13g2_decap_8
XFILLER_49_126 VDD VSS sg13g2_decap_8
XFILLER_92_405 VDD VSS sg13g2_fill_1
XFILLER_77_468 VDD VSS sg13g2_decap_8
XFILLER_73_630 VDD VSS sg13g2_decap_4
XFILLER_58_693 VDD VSS sg13g2_decap_8
XFILLER_38_84 VDD VSS sg13g2_decap_8
XFILLER_46_866 VDD VSS sg13g2_decap_8
XFILLER_18_546 VDD VSS sg13g2_decap_8
XFILLER_45_343 VDD VSS sg13g2_decap_8
XFILLER_61_858 VDD VSS sg13g2_decap_8
XFILLER_14_763 VDD VSS sg13g2_decap_8
XFILLER_13_273 VDD VSS sg13g2_decap_8
XFILLER_9_266 VDD VSS sg13g2_decap_8
Xclkload14 clkload14/Y _2345_/CLK VDD VSS sg13g2_inv_2
XFILLER_10_980 VDD VSS sg13g2_decap_8
XFILLER_86_1003 VDD VSS sg13g2_fill_2
XFILLER_6_973 VDD VSS sg13g2_decap_8
XFILLER_5_483 VDD VSS sg13g2_decap_8
X_1422_ _1422_/Y _1422_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_69_936 VDD VSS sg13g2_decap_8
XFILLER_96_700 VDD VSS sg13g2_decap_8
XFILLER_79_91 VDD VSS sg13g2_decap_8
XFILLER_68_413 VDD VSS sg13g2_decap_8
XFILLER_110_543 VDD VSS sg13g2_decap_8
XFILLER_84_906 VDD VSS sg13g2_decap_8
X_1353_ VDD _2205_/D _1353_/A VSS sg13g2_inv_1
XFILLER_84_917 VDD VSS sg13g2_fill_1
XFILLER_95_265 VDD VSS sg13g2_decap_8
X_1284_ _1284_/Y _1344_/B1 hold336/X _1344_/A2 _2336_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_1012 VDD VSS sg13g2_decap_8
XFILLER_83_438 VDD VSS sg13g2_decap_8
XFILLER_37_833 VDD VSS sg13g2_decap_8
XFILLER_76_490 VDD VSS sg13g2_fill_1
XFILLER_64_641 VDD VSS sg13g2_decap_8
XFILLER_36_343 VDD VSS sg13g2_decap_8
XFILLER_93_1018 VDD VSS sg13g2_decap_8
XFILLER_91_482 VDD VSS sg13g2_decap_8
XFILLER_63_173 VDD VSS sg13g2_fill_1
X_2176__188 VDD VSS _2176_/RESET_B sg13g2_tiehi
XFILLER_32_560 VDD VSS sg13g2_decap_8
XFILLER_51_368 VDD VSS sg13g2_decap_4
XFILLER_20_700 VDD VSS sg13g2_decap_8
Xclkload8 clkload8/Y clkload8/A VDD VSS sg13g2_inv_2
XFILLER_20_777 VDD VSS sg13g2_decap_8
XFILLER_30_1057 VDD VSS sg13g2_decap_4
XFILLER_105_337 VDD VSS sg13g2_decap_8
XFILLER_59_28 VDD VSS sg13g2_fill_2
XFILLER_8_1036 VDD VSS sg13g2_decap_8
XFILLER_87_766 VDD VSS sg13g2_decap_8
XFILLER_86_265 VDD VSS sg13g2_decap_4
XFILLER_59_457 VDD VSS sg13g2_decap_4
XFILLER_101_587 VDD VSS sg13g2_decap_8
XFILLER_74_438 VDD VSS sg13g2_decap_4
XFILLER_75_49 VDD VSS sg13g2_decap_8
XFILLER_28_833 VDD VSS sg13g2_decap_8
XFILLER_90_909 VDD VSS sg13g2_decap_8
XFILLER_55_641 VDD VSS sg13g2_decap_8
XFILLER_67_490 VDD VSS sg13g2_decap_8
XFILLER_27_343 VDD VSS sg13g2_decap_8
XFILLER_82_471 VDD VSS sg13g2_decap_8
XFILLER_43_814 VDD VSS sg13g2_decap_8
XFILLER_70_633 VDD VSS sg13g2_decap_8
XFILLER_39_1060 VDD VSS sg13g2_fill_1
XFILLER_23_560 VDD VSS sg13g2_decap_8
XFILLER_11_700 VDD VSS sg13g2_decap_8
XFILLER_24_42 VDD VSS sg13g2_decap_8
XFILLER_42_357 VDD VSS sg13g2_fill_2
XFILLER_10_210 VDD VSS sg13g2_decap_8
XFILLER_6_203 VDD VSS sg13g2_decap_8
XFILLER_11_777 VDD VSS sg13g2_decap_8
XFILLER_109_665 VDD VSS sg13g2_decap_8
XFILLER_10_287 VDD VSS sg13g2_decap_8
XFILLER_40_63 VDD VSS sg13g2_decap_8
XFILLER_108_175 VDD VSS sg13g2_decap_4
XFILLER_3_910 VDD VSS sg13g2_decap_8
XFILLER_2_420 VDD VSS sg13g2_decap_8
XFILLER_6_0 VDD VSS sg13g2_decap_8
XFILLER_112_819 VDD VSS sg13g2_decap_8
XFILLER_105_882 VDD VSS sg13g2_decap_8
XFILLER_78_711 VDD VSS sg13g2_decap_8
XFILLER_46_1031 VDD VSS sg13g2_decap_8
XFILLER_3_987 VDD VSS sg13g2_decap_8
XFILLER_111_329 VDD VSS sg13g2_decap_8
XFILLER_104_370 VDD VSS sg13g2_decap_8
XFILLER_77_221 VDD VSS sg13g2_decap_8
XFILLER_77_210 VDD VSS sg13g2_decap_8
XFILLER_2_497 VDD VSS sg13g2_decap_8
XFILLER_66_928 VDD VSS sg13g2_decap_8
XFILLER_77_287 VDD VSS sg13g2_decap_8
XFILLER_1_35 VDD VSS sg13g2_decap_8
XFILLER_19_833 VDD VSS sg13g2_decap_8
XFILLER_74_961 VDD VSS sg13g2_decap_8
XFILLER_92_235 VDD VSS sg13g2_decap_8
XFILLER_46_652 VDD VSS sg13g2_fill_2
XFILLER_58_490 VDD VSS sg13g2_decap_8
XFILLER_18_343 VDD VSS sg13g2_decap_8
XFILLER_61_611 VDD VSS sg13g2_decap_8
XFILLER_46_696 VDD VSS sg13g2_decap_8
XFILLER_34_847 VDD VSS sg13g2_decap_8
XFILLER_61_688 VDD VSS sg13g2_decap_8
XFILLER_61_666 VDD VSS sg13g2_decap_4
XFILLER_60_154 VDD VSS sg13g2_decap_8
XFILLER_33_357 VDD VSS sg13g2_decap_8
X_1971_ _1971_/B _1971_/C _1971_/A _2007_/B VDD VSS sg13g2_nand3_1
XFILLER_81_70 VDD VSS sg13g2_decap_8
XFILLER_14_560 VDD VSS sg13g2_decap_8
XFILLER_14_1008 VDD VSS sg13g2_decap_8
XFILLER_6_770 VDD VSS sg13g2_decap_8
XFILLER_5_280 VDD VSS sg13g2_decap_8
XFILLER_69_755 VDD VSS sg13g2_decap_8
X_1405_ _1406_/A _1392_/Y hold495/X _1392_/B _1385_/A VDD VSS sg13g2_a22oi_1
XFILLER_39_0 VDD VSS sg13g2_decap_8
X_1336_ _1336_/Y _1338_/B1 hold368/X _1338_/A2 _2331_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_340 VDD VSS sg13g2_decap_8
XFILLER_60_1039 VDD VSS sg13g2_decap_8
XFILLER_68_232 VDD VSS sg13g2_decap_8
XFILLER_56_405 VDD VSS sg13g2_decap_8
XFILLER_111_896 VDD VSS sg13g2_decap_8
XFILLER_96_585 VDD VSS sg13g2_decap_8
XFILLER_68_298 VDD VSS sg13g2_decap_8
X_1267_ VDD _2163_/D _1267_/A VSS sg13g2_inv_1
XFILLER_37_630 VDD VSS sg13g2_decap_8
XFILLER_65_972 VDD VSS sg13g2_decap_8
XFILLER_36_140 VDD VSS sg13g2_decap_8
X_1198_ VDD _1198_/Y _1198_/A VSS sg13g2_inv_1
XFILLER_92_791 VDD VSS sg13g2_decap_8
XFILLER_101_14 VDD VSS sg13g2_decap_8
XFILLER_25_847 VDD VSS sg13g2_decap_8
XFILLER_64_493 VDD VSS sg13g2_decap_8
XFILLER_52_677 VDD VSS sg13g2_decap_8
XFILLER_24_357 VDD VSS sg13g2_decap_8
X_2334__173 VDD VSS _2334_/RESET_B sg13g2_tiehi
XFILLER_20_574 VDD VSS sg13g2_decap_8
XFILLER_4_707 VDD VSS sg13g2_decap_8
XFILLER_69_1020 VDD VSS sg13g2_fill_1
X_2265__223 VDD VSS _2265_/RESET_B sg13g2_tiehi
XFILLER_3_217 VDD VSS sg13g2_decap_8
XFILLER_106_657 VDD VSS sg13g2_decap_8
XFILLER_105_112 VDD VSS sg13g2_decap_8
XFILLER_79_519 VDD VSS sg13g2_decap_8
XFILLER_10_77 VDD VSS sg13g2_decap_8
XFILLER_0_924 VDD VSS sg13g2_decap_8
XFILLER_102_874 VDD VSS sg13g2_decap_8
XFILLER_87_541 VDD VSS sg13g2_decap_8
XFILLER_59_243 VDD VSS sg13g2_decap_8
XFILLER_75_714 VDD VSS sg13g2_decap_8
XFILLER_101_351 VDD VSS sg13g2_decap_8
XFILLER_74_202 VDD VSS sg13g2_decap_8
XFILLER_59_298 VDD VSS sg13g2_fill_2
XFILLER_19_42 VDD VSS sg13g2_decap_8
XFILLER_63_909 VDD VSS sg13g2_decap_4
XFILLER_28_630 VDD VSS sg13g2_decap_8
XFILLER_90_717 VDD VSS sg13g2_decap_8
XFILLER_83_780 VDD VSS sg13g2_decap_8
XFILLER_74_279 VDD VSS sg13g2_decap_8
XFILLER_43_611 VDD VSS sg13g2_decap_8
XFILLER_27_140 VDD VSS sg13g2_decap_8
XFILLER_71_942 VDD VSS sg13g2_decap_8
XFILLER_16_847 VDD VSS sg13g2_decap_8
XFILLER_70_463 VDD VSS sg13g2_decap_8
XFILLER_37_1008 VDD VSS sg13g2_decap_8
XFILLER_15_357 VDD VSS sg13g2_decap_8
XFILLER_35_63 VDD VSS sg13g2_decap_8
XFILLER_43_688 VDD VSS sg13g2_decap_8
XFILLER_42_198 VDD VSS sg13g2_decap_8
XFILLER_11_574 VDD VSS sg13g2_decap_8
XFILLER_7_567 VDD VSS sg13g2_decap_8
XFILLER_51_95 VDD VSS sg13g2_fill_2
XFILLER_100_1011 VDD VSS sg13g2_decap_8
XFILLER_109_462 VDD VSS sg13g2_decap_8
XFILLER_83_1017 VDD VSS sg13g2_decap_8
XFILLER_98_806 VDD VSS sg13g2_decap_8
XFILLER_112_616 VDD VSS sg13g2_decap_8
XFILLER_111_126 VDD VSS sg13g2_decap_8
XFILLER_3_784 VDD VSS sg13g2_decap_8
XFILLER_32_7 VDD VSS sg13g2_decap_8
XFILLER_39_906 VDD VSS sg13g2_decap_8
XFILLER_2_294 VDD VSS sg13g2_decap_8
X_2170_ _2170_/RESET_B VSS VDD _2170_/D _2170_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_78_596 VDD VSS sg13g2_fill_2
XFILLER_78_585 VDD VSS sg13g2_decap_8
XFILLER_76_70 VDD VSS sg13g2_decap_8
XFILLER_66_714 VDD VSS sg13g2_decap_4
XFILLER_93_544 VDD VSS sg13g2_decap_4
XFILLER_47_950 VDD VSS sg13g2_decap_8
XFILLER_19_630 VDD VSS sg13g2_decap_8
XFILLER_20_1001 VDD VSS sg13g2_decap_8
XFILLER_18_140 VDD VSS sg13g2_decap_8
XFILLER_46_460 VDD VSS sg13g2_decap_4
XFILLER_80_227 VDD VSS sg13g2_decap_8
XFILLER_62_953 VDD VSS sg13g2_decap_8
XFILLER_34_644 VDD VSS sg13g2_decap_8
XFILLER_46_482 VDD VSS sg13g2_decap_8
XFILLER_33_154 VDD VSS sg13g2_decap_8
XFILLER_92_91 VDD VSS sg13g2_decap_8
XFILLER_61_474 VDD VSS sg13g2_decap_8
X_1954_ _1952_/A _1953_/Y _1954_/S _1955_/B VDD VSS sg13g2_mux2_1
XFILLER_30_861 VDD VSS sg13g2_decap_8
X_1885_ _1971_/B _1972_/A _1972_/B VDD VSS sg13g2_nand2_1
XFILLER_103_616 VDD VSS sg13g2_decap_8
XFILLER_89_817 VDD VSS sg13g2_decap_8
XFILLER_102_126 VDD VSS sg13g2_decap_8
XFILLER_96_371 VDD VSS sg13g2_decap_8
X_2368_ _2368_/RESET_B VSS VDD _2368_/D _2368_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_29_427 VDD VSS sg13g2_decap_8
XFILLER_111_693 VDD VSS sg13g2_decap_8
X_1319_ VDD _2189_/D _1319_/A VSS sg13g2_inv_1
XFILLER_84_544 VDD VSS sg13g2_decap_4
X_2299_ _2299_/RESET_B VSS VDD _2299_/D _2299_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_57_758 VDD VSS sg13g2_decap_8
XFILLER_56_235 VDD VSS sg13g2_decap_8
XFILLER_84_599 VDD VSS sg13g2_fill_2
XFILLER_72_717 VDD VSS sg13g2_decap_8
XFILLER_71_205 VDD VSS sg13g2_decap_8
XFILLER_38_961 VDD VSS sg13g2_decap_8
XFILLER_71_249 VDD VSS sg13g2_decap_8
XFILLER_112_35 VDD VSS sg13g2_decap_8
XFILLER_65_780 VDD VSS sg13g2_decap_8
XFILLER_25_644 VDD VSS sg13g2_decap_8
XFILLER_72_28 VDD VSS sg13g2_decap_8
XFILLER_52_452 VDD VSS sg13g2_fill_2
XFILLER_53_997 VDD VSS sg13g2_decap_8
XFILLER_24_154 VDD VSS sg13g2_decap_8
XFILLER_40_669 VDD VSS sg13g2_decap_8
XFILLER_21_861 VDD VSS sg13g2_decap_8
XFILLER_20_371 VDD VSS sg13g2_decap_8
XFILLER_21_21 VDD VSS sg13g2_decap_8
XFILLER_107_933 VDD VSS sg13g2_decap_8
XFILLER_4_504 VDD VSS sg13g2_decap_8
XFILLER_106_421 VDD VSS sg13g2_decap_8
XFILLER_97_14 VDD VSS sg13g2_decap_8
XFILLER_21_98 VDD VSS sg13g2_decap_8
XIO_BOND_vdd_pads\[0\].vdd_pad VDD bondpad_70x70
XFILLER_79_327 VDD VSS sg13g2_decap_8
XFILLER_0_721 VDD VSS sg13g2_decap_8
XFILLER_88_872 VDD VSS sg13g2_decap_8
XFILLER_75_500 VDD VSS sg13g2_decap_4
XFILLER_43_1045 VDD VSS sg13g2_decap_8
XFILLER_0_798 VDD VSS sg13g2_decap_8
XFILLER_102_693 VDD VSS sg13g2_decap_8
XFILLER_47_224 VDD VSS sg13g2_decap_8
XFILLER_75_588 VDD VSS sg13g2_decap_8
XFILLER_47_257 VDD VSS sg13g2_decap_8
XFILLER_44_942 VDD VSS sg13g2_decap_8
XFILLER_29_994 VDD VSS sg13g2_decap_8
XFILLER_56_791 VDD VSS sg13g2_decap_8
XFILLER_62_216 VDD VSS sg13g2_fill_2
XFILLER_46_84 VDD VSS sg13g2_decap_8
XFILLER_16_644 VDD VSS sg13g2_decap_8
XFILLER_43_441 VDD VSS sg13g2_decap_8
XFILLER_15_154 VDD VSS sg13g2_decap_8
XFILLER_31_658 VDD VSS sg13g2_decap_8
XFILLER_12_861 VDD VSS sg13g2_decap_8
XFILLER_30_168 VDD VSS sg13g2_decap_8
XFILLER_50_1038 VDD VSS sg13g2_decap_8
XFILLER_11_371 VDD VSS sg13g2_decap_8
XFILLER_8_854 VDD VSS sg13g2_decap_8
X_1670_ _1670_/A _1670_/B _2306_/D VDD VSS sg13g2_nor2_1
XFILLER_7_364 VDD VSS sg13g2_decap_8
XFILLER_7_56 VDD VSS sg13g2_decap_8
Xhold309 _1300_/Y VDD VSS _1301_/A sg13g2_dlygate4sd3_1
X_2248__251 VDD VSS _2248_/RESET_B sg13g2_tiehi
XFILLER_112_413 VDD VSS sg13g2_decap_8
XFILLER_3_581 VDD VSS sg13g2_decap_8
XFILLER_86_809 VDD VSS sg13g2_decap_8
XFILLER_97_179 VDD VSS sg13g2_decap_8
X_2222_ _2222__96/L_HI VSS VDD _2222_/D _2222_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_87_91 VDD VSS sg13g2_decap_8
XFILLER_39_703 VDD VSS sg13g2_decap_8
X_2153_ _2162_/B _2040_/A _2332_/D VDD VSS sg13g2_nor2b_1
XFILLER_93_330 VDD VSS sg13g2_fill_2
XFILLER_78_382 VDD VSS sg13g2_decap_8
XFILLER_66_533 VDD VSS sg13g2_decap_8
XFILLER_38_224 VDD VSS sg13g2_decap_8
XFILLER_93_341 VDD VSS sg13g2_decap_8
XFILLER_81_503 VDD VSS sg13g2_decap_8
XFILLER_54_728 VDD VSS sg13g2_decap_8
XFILLER_4_1050 VDD VSS sg13g2_decap_8
X_2084_ _2080_/Y VDD _2341_/D VSS _2082_/Y _2083_/Y sg13g2_o21ai_1
XFILLER_35_931 VDD VSS sg13g2_decap_8
XFILLER_66_599 VDD VSS sg13g2_decap_8
XFILLER_53_238 VDD VSS sg13g2_decap_8
XFILLER_59_1041 VDD VSS sg13g2_decap_8
XFILLER_62_761 VDD VSS sg13g2_decap_8
XFILLER_34_441 VDD VSS sg13g2_decap_8
XFILLER_62_794 VDD VSS sg13g2_fill_1
XFILLER_107_1017 VDD VSS sg13g2_decap_8
XFILLER_50_967 VDD VSS sg13g2_decap_8
XFILLER_22_658 VDD VSS sg13g2_decap_8
XFILLER_21_168 VDD VSS sg13g2_decap_8
X_1937_ _1935_/Y _1936_/Y _1954_/S _1938_/B VDD VSS sg13g2_mux2_1
X_1868_ _1866_/A _1854_/A _1854_/C _1869_/B VDD VSS sg13g2_a21o_1
X_1799_ _1825_/A _1823_/A _1800_/C VDD VSS sg13g2_nor2_1
XFILLER_104_936 VDD VSS sg13g2_decap_8
XFILLER_103_413 VDD VSS sg13g2_fill_2
XFILLER_107_35 VDD VSS sg13g2_decap_8
XFILLER_66_1056 VDD VSS sg13g2_decap_4
XFILLER_1_518 VDD VSS sg13g2_decap_8
XFILLER_77_809 VDD VSS sg13g2_decap_8
XFILLER_27_1029 VDD VSS sg13g2_decap_8
XFILLER_67_28 VDD VSS sg13g2_decap_8
XFILLER_112_980 VDD VSS sg13g2_decap_8
XFILLER_88_168 VDD VSS sg13g2_fill_2
XFILLER_57_500 VDD VSS sg13g2_decap_8
XFILLER_85_831 VDD VSS sg13g2_decap_4
XFILLER_111_490 VDD VSS sg13g2_decap_8
XFILLER_69_393 VDD VSS sg13g2_decap_8
XFILLER_29_224 VDD VSS sg13g2_decap_8
XFILLER_84_341 VDD VSS sg13g2_decap_8
XFILLER_57_588 VDD VSS sg13g2_fill_2
XFILLER_84_385 VDD VSS sg13g2_decap_8
XFILLER_72_536 VDD VSS sg13g2_decap_8
XFILLER_83_49 VDD VSS sg13g2_decap_8
XFILLER_26_931 VDD VSS sg13g2_decap_8
XFILLER_44_227 VDD VSS sg13g2_fill_1
XFILLER_16_21 VDD VSS sg13g2_decap_8
XFILLER_25_441 VDD VSS sg13g2_decap_8
XFILLER_73_1016 VDD VSS sg13g2_decap_8
XFILLER_41_923 VDD VSS sg13g2_decap_8
XFILLER_80_591 VDD VSS sg13g2_decap_8
XFILLER_16_98 VDD VSS sg13g2_decap_8
XFILLER_13_658 VDD VSS sg13g2_decap_8
XFILLER_40_433 VDD VSS sg13g2_decap_8
XFILLER_52_293 VDD VSS sg13g2_decap_8
XFILLER_12_168 VDD VSS sg13g2_decap_8
XFILLER_40_477 VDD VSS sg13g2_decap_8
XFILLER_32_42 VDD VSS sg13g2_decap_8
XFILLER_107_730 VDD VSS sg13g2_decap_8
XFILLER_4_301 VDD VSS sg13g2_decap_8
XFILLER_10_1022 VDD VSS sg13g2_decap_8
XFILLER_106_0 VDD VSS sg13g2_decap_8
XFILLER_5_868 VDD VSS sg13g2_decap_8
XFILLER_106_273 VDD VSS sg13g2_decap_8
XFILLER_4_378 VDD VSS sg13g2_decap_8
XFILLER_110_928 VDD VSS sg13g2_decap_8
XFILLER_103_980 VDD VSS sg13g2_decap_8
X_2204__132 VDD VSS _2204_/RESET_B sg13g2_tiehi
XFILLER_94_105 VDD VSS sg13g2_decap_8
XFILLER_67_308 VDD VSS sg13g2_decap_8
XFILLER_87_190 VDD VSS sg13g2_decap_8
XFILLER_0_595 VDD VSS sg13g2_decap_8
XFILLER_91_801 VDD VSS sg13g2_decap_8
XFILLER_76_886 VDD VSS sg13g2_decap_8
XFILLER_75_341 VDD VSS sg13g2_decap_8
XFILLER_36_728 VDD VSS sg13g2_decap_8
XFILLER_29_791 VDD VSS sg13g2_decap_8
XFILLER_17_931 VDD VSS sg13g2_decap_8
XFILLER_35_238 VDD VSS sg13g2_decap_8
XFILLER_90_333 VDD VSS sg13g2_decap_8
XFILLER_16_441 VDD VSS sg13g2_decap_8
XFILLER_71_591 VDD VSS sg13g2_decap_8
XFILLER_32_945 VDD VSS sg13g2_decap_8
XFILLER_31_455 VDD VSS sg13g2_decap_8
X_1722_ _1725_/A _1722_/B _1722_/Y VDD VSS sg13g2_nor2_1
XFILLER_8_651 VDD VSS sg13g2_decap_8
X_1653_ _1674_/B _2330_/Q _2322_/Q _2345_/Q _2337_/Q _1677_/A _1653_/X VDD VSS sg13g2_mux4_1
XFILLER_7_161 VDD VSS sg13g2_decap_8
XFILLER_99_945 VDD VSS sg13g2_decap_8
XFILLER_112_210 VDD VSS sg13g2_decap_8
XFILLER_98_411 VDD VSS sg13g2_decap_8
X_1584_ _2285_/D _1589_/C _1584_/B _2284_/D VDD VSS sg13g2_and3_1
XIO_FILL_IO_EAST_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_85_105 VDD VSS sg13g2_decap_8
XFILLER_67_820 VDD VSS sg13g2_decap_8
XFILLER_21_0 VDD VSS sg13g2_decap_8
XFILLER_112_287 VDD VSS sg13g2_decap_8
X_2205_ _2205_/RESET_B VSS VDD _2205_/D _2205_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_522 VDD VSS sg13g2_fill_1
XFILLER_39_577 VDD VSS sg13g2_decap_8
X_2136_ _2124_/A _2200_/Q _2192_/Q _2184_/Q _2176_/Q _2144_/S1 _2136_/X VDD VSS sg13g2_mux4_1
XFILLER_94_683 VDD VSS sg13g2_decap_4
XFILLER_82_834 VDD VSS sg13g2_decap_8
XFILLER_93_171 VDD VSS sg13g2_decap_8
XFILLER_27_728 VDD VSS sg13g2_decap_8
XFILLER_66_385 VDD VSS sg13g2_decap_8
XFILLER_54_536 VDD VSS sg13g2_fill_1
X_2067_ _2055_/B _2056_/X _2079_/S _2068_/B VDD VSS sg13g2_mux2_1
XFILLER_81_333 VDD VSS sg13g2_decap_8
XFILLER_26_238 VDD VSS sg13g2_decap_8
XFILLER_23_945 VDD VSS sg13g2_decap_8
XFILLER_50_742 VDD VSS sg13g2_decap_8
XFILLER_72_1060 VDD VSS sg13g2_fill_1
XFILLER_22_455 VDD VSS sg13g2_decap_8
XFILLER_33_1022 VDD VSS sg13g2_decap_8
XFILLER_108_549 VDD VSS sg13g2_decap_8
X_2186__168 VDD VSS _2186_/RESET_B sg13g2_tiehi
XFILLER_2_805 VDD VSS sg13g2_decap_8
XFILLER_104_722 VDD VSS sg13g2_decap_8
XFILLER_78_49 VDD VSS sg13g2_decap_8
XFILLER_1_315 VDD VSS sg13g2_decap_8
XFILLER_89_444 VDD VSS sg13g2_decap_8
XFILLER_89_433 VDD VSS sg13g2_decap_8
XFILLER_104_799 VDD VSS sg13g2_decap_8
XFILLER_77_639 VDD VSS sg13g2_decap_8
XFILLER_76_105 VDD VSS sg13g2_decap_8
XFILLER_85_661 VDD VSS sg13g2_decap_8
XFILLER_40_1026 VDD VSS sg13g2_decap_8
XFILLER_57_330 VDD VSS sg13g2_decap_8
XFILLER_100_994 VDD VSS sg13g2_decap_4
XFILLER_18_728 VDD VSS sg13g2_decap_8
XFILLER_27_42 VDD VSS sg13g2_decap_8
XFILLER_45_525 VDD VSS sg13g2_decap_8
XFILLER_17_238 VDD VSS sg13g2_decap_8
XFILLER_72_366 VDD VSS sg13g2_decap_8
XFILLER_60_517 VDD VSS sg13g2_decap_8
XFILLER_53_580 VDD VSS sg13g2_decap_8
XFILLER_41_720 VDD VSS sg13g2_decap_8
XFILLER_14_945 VDD VSS sg13g2_decap_8
XFILLER_13_455 VDD VSS sg13g2_decap_8
XFILLER_43_63 VDD VSS sg13g2_decap_8
XFILLER_40_252 VDD VSS sg13g2_decap_8
XFILLER_41_797 VDD VSS sg13g2_decap_8
XFILLER_9_448 VDD VSS sg13g2_decap_8
XFILLER_5_665 VDD VSS sg13g2_decap_8
XFILLER_4_175 VDD VSS sg13g2_decap_8
X_2245__254 VDD VSS _2245_/RESET_B sg13g2_tiehi
XFILLER_4_35 VDD VSS sg13g2_decap_8
XFILLER_110_725 VDD VSS sg13g2_decap_8
XFILLER_67_105 VDD VSS sg13g2_decap_8
XFILLER_68_60 VDD VSS sg13g2_fill_1
XFILLER_68_71 VDD VSS sg13g2_fill_1
XFILLER_1_882 VDD VSS sg13g2_decap_8
XFILLER_68_82 VDD VSS sg13g2_decap_8
XFILLER_76_650 VDD VSS sg13g2_decap_8
XFILLER_95_469 VDD VSS sg13g2_decap_8
XFILLER_0_392 VDD VSS sg13g2_decap_8
XFILLER_75_171 VDD VSS sg13g2_decap_8
XFILLER_64_823 VDD VSS sg13g2_decap_8
XFILLER_49_897 VDD VSS sg13g2_decap_8
XFILLER_63_311 VDD VSS sg13g2_decap_8
XFILLER_36_525 VDD VSS sg13g2_decap_8
XFILLER_48_374 VDD VSS sg13g2_decap_8
XFILLER_84_70 VDD VSS sg13g2_decap_8
XFILLER_91_697 VDD VSS sg13g2_decap_8
XFILLER_90_174 VDD VSS sg13g2_decap_8
XFILLER_63_366 VDD VSS sg13g2_decap_8
XFILLER_56_1022 VDD VSS sg13g2_decap_8
XFILLER_32_742 VDD VSS sg13g2_decap_8
X_2252__247 VDD VSS _2252_/RESET_B sg13g2_tiehi
XFILLER_31_252 VDD VSS sg13g2_decap_8
XFILLER_20_959 VDD VSS sg13g2_decap_8
X_1705_ _1705_/Y _1720_/A _1705_/B VDD VSS sg13g2_nand2_1
XFILLER_69_0 VDD VSS sg13g2_decap_8
XFILLER_105_519 VDD VSS sg13g2_decap_8
X_1636_ _1639_/A _1636_/B _1636_/Y VDD VSS sg13g2_nor2_1
X_1567_ _1566_/Y VDD _1567_/Y VSS _2288_/Q _1564_/Y sg13g2_o21ai_1
XFILLER_98_274 VDD VSS sg13g2_decap_8
XFILLER_101_758 VDD VSS sg13g2_decap_8
XFILLER_100_202 VDD VSS sg13g2_fill_2
XFILLER_86_447 VDD VSS sg13g2_decap_8
X_1498_ _1236_/C VDD _1498_/Y VSS hold295/X _1497_/B sg13g2_o21ai_1
XFILLER_100_268 VDD VSS sg13g2_decap_8
XFILLER_104_14 VDD VSS sg13g2_decap_8
XFILLER_58_149 VDD VSS sg13g2_decap_8
XFILLER_39_352 VDD VSS sg13g2_decap_8
XFILLER_73_119 VDD VSS sg13g2_decap_8
XFILLER_66_160 VDD VSS sg13g2_decap_8
XFILLER_27_525 VDD VSS sg13g2_decap_8
XFILLER_82_653 VDD VSS sg13g2_decap_8
X_2119_ VSS VDD _2144_/S0 _1218_/Y _2120_/B _2118_/Y sg13g2_a21oi_1
XFILLER_55_867 VDD VSS sg13g2_decap_8
XFILLER_70_815 VDD VSS sg13g2_decap_8
XFILLER_54_366 VDD VSS sg13g2_decap_8
Xfanout12 _1990_/Y _2036_/S VDD VSS sg13g2_buf_1
XFILLER_23_742 VDD VSS sg13g2_decap_8
Xfanout45 _2356_/Q _2142_/A1 VDD VSS sg13g2_buf_1
XFILLER_80_28 VDD VSS sg13g2_decap_8
Xfanout34 _1342_/A2 _1482_/A2 VDD VSS sg13g2_buf_1
Xfanout23 _1481_/A2 _1479_/A2 VDD VSS sg13g2_buf_1
XFILLER_22_252 VDD VSS sg13g2_decap_8
Xfanout56 _2286_/Q _1577_/S0 VDD VSS sg13g2_buf_1
Xfanout67 _2106_/A _2101_/A VDD VSS sg13g2_buf_1
Xfanout78 fanout78/A _2138_/B1 VDD VSS sg13g2_buf_1
XFILLER_11_959 VDD VSS sg13g2_decap_8
XFILLER_10_469 VDD VSS sg13g2_decap_8
XFILLER_109_847 VDD VSS sg13g2_decap_8
XFILLER_13_77 VDD VSS sg13g2_decap_8
XFILLER_2_602 VDD VSS sg13g2_decap_8
XFILLER_89_230 VDD VSS sg13g2_decap_8
Xhold481 _2212_/Q VDD VSS _1371_/A sg13g2_dlygate4sd3_1
Xhold470 _2205_/Q VDD VSS hold470/X sg13g2_dlygate4sd3_1
XFILLER_1_112 VDD VSS sg13g2_decap_8
XFILLER_78_937 VDD VSS sg13g2_decap_8
XFILLER_104_563 VDD VSS sg13g2_decap_8
Xhold492 _1690_/Y VDD VSS _2313_/D sg13g2_dlygate4sd3_1
XFILLER_2_679 VDD VSS sg13g2_decap_8
XFILLER_77_436 VDD VSS sg13g2_decap_8
XFILLER_1_189 VDD VSS sg13g2_decap_8
XFILLER_38_63 VDD VSS sg13g2_decap_8
XFILLER_58_672 VDD VSS sg13g2_decap_8
X_2275__203 VDD VSS _2275_/RESET_B sg13g2_tiehi
XFILLER_18_525 VDD VSS sg13g2_decap_8
XFILLER_73_653 VDD VSS sg13g2_decap_8
XFILLER_46_856 VDD VSS sg13g2_fill_1
XFILLER_57_193 VDD VSS sg13g2_decap_8
XFILLER_45_322 VDD VSS sg13g2_decap_8
XFILLER_45_388 VDD VSS sg13g2_decap_8
XFILLER_72_196 VDD VSS sg13g2_decap_8
XFILLER_14_742 VDD VSS sg13g2_decap_8
XFILLER_33_539 VDD VSS sg13g2_decap_8
XFILLER_41_550 VDD VSS sg13g2_decap_8
XFILLER_13_252 VDD VSS sg13g2_decap_8
XFILLER_41_594 VDD VSS sg13g2_decap_8
XFILLER_9_245 VDD VSS sg13g2_decap_8
XFILLER_16_1050 VDD VSS sg13g2_decap_8
Xclkload15 _2337_/CLK clkload15/Y VDD VSS sg13g2_inv_4
XFILLER_6_952 VDD VSS sg13g2_decap_8
XFILLER_62_7 VDD VSS sg13g2_decap_8
XFILLER_86_1059 VDD VSS sg13g2_fill_2
XFILLER_86_1048 VDD VSS sg13g2_decap_8
XFILLER_5_462 VDD VSS sg13g2_decap_8
X_1421_ _1420_/Y VDD _2231_/D VSS _1379_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_79_70 VDD VSS sg13g2_decap_8
XFILLER_69_915 VDD VSS sg13g2_decap_8
XFILLER_110_522 VDD VSS sg13g2_decap_8
X_1352_ _1353_/A _1347_/Y hold470/X _1347_/B _1373_/A VDD VSS sg13g2_a22oi_1
XFILLER_96_789 VDD VSS sg13g2_decap_8
XFILLER_95_255 VDD VSS sg13g2_fill_2
X_1283_ VDD _2171_/D _1283_/A VSS sg13g2_inv_1
XFILLER_56_609 VDD VSS sg13g2_decap_8
XFILLER_110_599 VDD VSS sg13g2_decap_8
XFILLER_83_417 VDD VSS sg13g2_decap_8
XFILLER_95_91 VDD VSS sg13g2_decap_8
XFILLER_23_1043 VDD VSS sg13g2_decap_8
XFILLER_64_620 VDD VSS sg13g2_decap_8
XFILLER_49_683 VDD VSS sg13g2_decap_8
XFILLER_37_812 VDD VSS sg13g2_decap_8
XFILLER_36_322 VDD VSS sg13g2_decap_8
XFILLER_48_182 VDD VSS sg13g2_decap_8
XFILLER_91_461 VDD VSS sg13g2_decap_8
XFILLER_37_889 VDD VSS sg13g2_decap_8
XFILLER_63_152 VDD VSS sg13g2_decap_8
XFILLER_64_697 VDD VSS sg13g2_decap_8
XFILLER_51_347 VDD VSS sg13g2_decap_8
XFILLER_24_539 VDD VSS sg13g2_decap_8
XFILLER_36_399 VDD VSS sg13g2_decap_8
Xclkload9 VDD clkload9/Y clkload9/A VSS sg13g2_inv_1
XFILLER_20_756 VDD VSS sg13g2_decap_8
XFILLER_30_1036 VDD VSS sg13g2_decap_8
XFILLER_106_839 VDD VSS sg13g2_decap_8
XFILLER_105_316 VDD VSS sg13g2_decap_8
X_1619_ _1619_/Y _1638_/S _1619_/B VDD VSS sg13g2_nand2_1
XFILLER_8_1015 VDD VSS sg13g2_decap_8
XFILLER_99_583 VDD VSS sg13g2_decap_8
XFILLER_87_745 VDD VSS sg13g2_decap_8
XFILLER_75_918 VDD VSS sg13g2_decap_8
XFILLER_101_566 VDD VSS sg13g2_decap_8
XFILLER_86_244 VDD VSS sg13g2_decap_8
XFILLER_75_28 VDD VSS sg13g2_decap_8
XFILLER_47_609 VDD VSS sg13g2_decap_8
XFILLER_86_299 VDD VSS sg13g2_decap_8
XFILLER_74_417 VDD VSS sg13g2_decap_8
XFILLER_55_620 VDD VSS sg13g2_decap_8
XFILLER_28_812 VDD VSS sg13g2_decap_8
XFILLER_27_322 VDD VSS sg13g2_decap_8
XFILLER_39_182 VDD VSS sg13g2_decap_8
XFILLER_70_612 VDD VSS sg13g2_decap_8
XFILLER_82_450 VDD VSS sg13g2_decap_4
XFILLER_28_889 VDD VSS sg13g2_decap_8
XFILLER_54_141 VDD VSS sg13g2_decap_8
XFILLER_91_49 VDD VSS sg13g2_decap_8
XFILLER_54_196 VDD VSS sg13g2_decap_8
XFILLER_15_539 VDD VSS sg13g2_decap_8
XFILLER_27_399 VDD VSS sg13g2_decap_8
XFILLER_42_325 VDD VSS sg13g2_fill_2
XFILLER_42_336 VDD VSS sg13g2_decap_8
XFILLER_70_689 VDD VSS sg13g2_decap_8
XFILLER_24_21 VDD VSS sg13g2_decap_8
XFILLER_11_756 VDD VSS sg13g2_decap_8
XFILLER_24_98 VDD VSS sg13g2_decap_8
XFILLER_10_266 VDD VSS sg13g2_decap_8
XFILLER_7_749 VDD VSS sg13g2_decap_8
XFILLER_109_644 VDD VSS sg13g2_decap_8
XFILLER_6_259 VDD VSS sg13g2_decap_8
XFILLER_40_42 VDD VSS sg13g2_decap_8
XFILLER_108_154 VDD VSS sg13g2_decap_8
XFILLER_105_861 VDD VSS sg13g2_decap_8
XFILLER_111_308 VDD VSS sg13g2_decap_8
XFILLER_46_1010 VDD VSS sg13g2_decap_8
XFILLER_3_966 VDD VSS sg13g2_decap_8
XFILLER_2_476 VDD VSS sg13g2_decap_8
XFILLER_78_789 VDD VSS sg13g2_decap_8
XFILLER_66_907 VDD VSS sg13g2_decap_8
XFILLER_1_14 VDD VSS sg13g2_decap_8
XFILLER_92_214 VDD VSS sg13g2_decap_8
XFILLER_77_266 VDD VSS sg13g2_decap_8
XFILLER_59_992 VDD VSS sg13g2_decap_8
XFILLER_65_406 VDD VSS sg13g2_decap_8
XFILLER_19_812 VDD VSS sg13g2_decap_8
XFILLER_37_119 VDD VSS sg13g2_decap_8
XFILLER_74_940 VDD VSS sg13g2_decap_8
XFILLER_93_759 VDD VSS sg13g2_decap_8
XFILLER_18_322 VDD VSS sg13g2_decap_8
XFILLER_73_450 VDD VSS sg13g2_fill_1
XFILLER_34_826 VDD VSS sg13g2_decap_8
XFILLER_19_889 VDD VSS sg13g2_decap_8
XFILLER_65_94 VDD VSS sg13g2_decap_8
XFILLER_61_645 VDD VSS sg13g2_fill_2
XFILLER_18_399 VDD VSS sg13g2_decap_8
XFILLER_33_336 VDD VSS sg13g2_decap_8
XFILLER_45_196 VDD VSS sg13g2_decap_8
X_1970_ _1973_/B _1973_/A _1886_/Y _1971_/C VDD VSS sg13g2_a21o_1
XFILLER_61_678 VDD VSS sg13g2_fill_1
XFILLER_61_656 VDD VSS sg13g2_decap_8
XFILLER_60_133 VDD VSS sg13g2_decap_8
XFILLER_53_1047 VDD VSS sg13g2_decap_8
XFILLER_69_734 VDD VSS sg13g2_decap_8
X_1404_ VDD _2224_/D _1404_/A VSS sg13g2_inv_1
XFILLER_102_319 VDD VSS sg13g2_decap_8
XFILLER_68_211 VDD VSS sg13g2_decap_8
XFILLER_111_875 VDD VSS sg13g2_decap_8
XFILLER_96_542 VDD VSS sg13g2_fill_1
XFILLER_96_564 VDD VSS sg13g2_decap_8
X_1335_ VDD _2197_/D _1335_/A VSS sg13g2_inv_1
XFILLER_60_1018 VDD VSS sg13g2_decap_8
XFILLER_57_929 VDD VSS sg13g2_decap_8
XFILLER_29_609 VDD VSS sg13g2_decap_8
XFILLER_84_726 VDD VSS sg13g2_decap_8
XFILLER_68_277 VDD VSS sg13g2_decap_8
XFILLER_28_119 VDD VSS sg13g2_decap_8
XFILLER_110_396 VDD VSS sg13g2_decap_8
XFILLER_83_247 VDD VSS sg13g2_fill_2
XFILLER_65_951 VDD VSS sg13g2_decap_8
X_1266_ _1266_/Y _1280_/B1 hold379/X _1280_/A2 _2313_/Q VDD VSS sg13g2_a22oi_1
XFILLER_92_770 VDD VSS sg13g2_decap_8
XFILLER_37_686 VDD VSS sg13g2_decap_8
XFILLER_25_826 VDD VSS sg13g2_decap_8
X_1197_ VDD _1197_/Y _1242_/B VSS sg13g2_inv_1
XFILLER_91_280 VDD VSS sg13g2_fill_2
XFILLER_52_645 VDD VSS sg13g2_decap_8
XFILLER_64_472 VDD VSS sg13g2_decap_8
XFILLER_24_336 VDD VSS sg13g2_decap_8
XFILLER_36_196 VDD VSS sg13g2_decap_8
XFILLER_80_987 VDD VSS sg13g2_decap_8
XFILLER_52_656 VDD VSS sg13g2_fill_1
XFILLER_51_133 VDD VSS sg13g2_decap_8
XFILLER_51_188 VDD VSS sg13g2_decap_8
X_2369__226 VDD VSS _2369_/RESET_B sg13g2_tiehi
XFILLER_20_553 VDD VSS sg13g2_decap_8
XFILLER_106_636 VDD VSS sg13g2_decap_8
XFILLER_10_56 VDD VSS sg13g2_decap_8
XFILLER_0_903 VDD VSS sg13g2_decap_8
XFILLER_99_380 VDD VSS sg13g2_decap_8
XFILLER_59_222 VDD VSS sg13g2_decap_8
XFILLER_102_853 VDD VSS sg13g2_decap_8
XFILLER_101_330 VDD VSS sg13g2_decap_8
XFILLER_86_49 VDD VSS sg13g2_decap_8
XFILLER_19_21 VDD VSS sg13g2_decap_8
XFILLER_87_597 VDD VSS sg13g2_decap_8
XFILLER_19_119 VDD VSS sg13g2_decap_8
XFILLER_47_406 VDD VSS sg13g2_fill_2
XFILLER_47_428 VDD VSS sg13g2_decap_8
XFILLER_19_98 VDD VSS sg13g2_decap_8
XFILLER_74_258 VDD VSS sg13g2_decap_8
XFILLER_56_984 VDD VSS sg13g2_decap_8
XFILLER_16_826 VDD VSS sg13g2_decap_8
XFILLER_71_921 VDD VSS sg13g2_decap_8
XFILLER_28_686 VDD VSS sg13g2_decap_8
XFILLER_55_494 VDD VSS sg13g2_decap_8
XFILLER_15_336 VDD VSS sg13g2_decap_8
XFILLER_35_42 VDD VSS sg13g2_decap_8
XFILLER_76_1058 VDD VSS sg13g2_fill_2
XFILLER_70_442 VDD VSS sg13g2_decap_8
XFILLER_70_431 VDD VSS sg13g2_fill_1
XIO_BOND_out_data_pads\[2\].out_data_pad out_data_PADs[2] bondpad_70x70
XFILLER_43_667 VDD VSS sg13g2_decap_8
XFILLER_42_133 VDD VSS sg13g2_decap_8
XFILLER_27_196 VDD VSS sg13g2_decap_8
XFILLER_71_998 VDD VSS sg13g2_decap_8
XFILLER_42_177 VDD VSS sg13g2_decap_8
XFILLER_11_553 VDD VSS sg13g2_decap_8
XFILLER_109_441 VDD VSS sg13g2_decap_8
XFILLER_7_546 VDD VSS sg13g2_decap_8
XFILLER_51_74 VDD VSS sg13g2_decap_8
XFILLER_3_763 VDD VSS sg13g2_decap_8
XFILLER_111_105 VDD VSS sg13g2_decap_8
XFILLER_2_273 VDD VSS sg13g2_decap_8
XFILLER_25_7 VDD VSS sg13g2_decap_8
XFILLER_93_512 VDD VSS sg13g2_decap_8
XFILLER_65_247 VDD VSS sg13g2_decap_8
XFILLER_38_439 VDD VSS sg13g2_decap_8
Xin_data_pads\[3\].in_data_pad IOVDD IOVSS _1376_/A in_data_PADs[3] VDD VSS sg13g2_IOPadIn
XFILLER_81_729 VDD VSS sg13g2_decap_8
XFILLER_80_206 VDD VSS sg13g2_decap_8
XFILLER_65_269 VDD VSS sg13g2_decap_8
XFILLER_62_921 VDD VSS sg13g2_fill_1
XFILLER_34_623 VDD VSS sg13g2_decap_8
XFILLER_19_686 VDD VSS sg13g2_decap_8
XFILLER_20_1057 VDD VSS sg13g2_decap_4
XFILLER_92_70 VDD VSS sg13g2_decap_8
XFILLER_61_453 VDD VSS sg13g2_decap_8
XFILLER_18_196 VDD VSS sg13g2_decap_8
XFILLER_33_133 VDD VSS sg13g2_decap_8
X_2214__112 VDD VSS _2214_/RESET_B sg13g2_tiehi
X_1953_ VDD _1953_/Y _1953_/A VSS sg13g2_inv_1
XFILLER_30_840 VDD VSS sg13g2_decap_8
X_1884_ _1972_/B _1884_/A _1884_/B VDD VSS sg13g2_xnor2_1
XIO_FILL_IO_SOUTH_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_51_0 VDD VSS sg13g2_decap_8
XFILLER_88_339 VDD VSS sg13g2_decap_8
XFILLER_102_105 VDD VSS sg13g2_decap_8
XFILLER_99_1014 VDD VSS sg13g2_decap_4
XFILLER_111_672 VDD VSS sg13g2_decap_8
XFILLER_97_895 VDD VSS sg13g2_decap_8
XFILLER_69_586 VDD VSS sg13g2_decap_8
XFILLER_96_350 VDD VSS sg13g2_decap_8
X_2367_ _2367_/RESET_B VSS VDD _2367_/D _2367_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_57_737 VDD VSS sg13g2_decap_8
XFILLER_5_1029 VDD VSS sg13g2_decap_8
XFILLER_29_406 VDD VSS sg13g2_decap_8
XFILLER_99_1025 VDD VSS sg13g2_fill_1
X_1318_ _1318_/Y _1322_/B1 hold377/X _1322_/A2 _2322_/Q VDD VSS sg13g2_a22oi_1
XFILLER_84_556 VDD VSS sg13g2_decap_8
XFILLER_110_182 VDD VSS sg13g2_decap_8
XFILLER_84_523 VDD VSS sg13g2_decap_8
XFILLER_38_940 VDD VSS sg13g2_decap_8
X_2298_ _2298_/RESET_B VSS VDD _2298_/D _2298_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_112_14 VDD VSS sg13g2_decap_8
X_1249_ _1249_/A _1249_/B _1249_/C _1250_/B VDD VSS sg13g2_nor3_1
XFILLER_65_792 VDD VSS sg13g2_decap_8
XFILLER_25_623 VDD VSS sg13g2_decap_8
XFILLER_37_483 VDD VSS sg13g2_decap_8
XFILLER_53_976 VDD VSS sg13g2_decap_8
XFILLER_52_431 VDD VSS sg13g2_decap_8
XFILLER_24_133 VDD VSS sg13g2_decap_8
XFILLER_40_648 VDD VSS sg13g2_decap_8
XFILLER_21_840 VDD VSS sg13g2_decap_8
XFILLER_20_350 VDD VSS sg13g2_decap_8
X_2232__289 VDD VSS _2232_/RESET_B sg13g2_tiehi
XFILLER_107_912 VDD VSS sg13g2_decap_8
XFILLER_106_400 VDD VSS sg13g2_decap_8
XFILLER_21_77 VDD VSS sg13g2_decap_8
XFILLER_107_989 VDD VSS sg13g2_decap_8
XFILLER_106_477 VDD VSS sg13g2_decap_8
XFILLER_106_488 VDD VSS sg13g2_fill_1
XFILLER_0_700 VDD VSS sg13g2_decap_8
XFILLER_82_1040 VDD VSS sg13g2_decap_8
XFILLER_88_851 VDD VSS sg13g2_decap_8
XFILLER_43_1024 VDD VSS sg13g2_decap_8
XFILLER_48_715 VDD VSS sg13g2_fill_2
XFILLER_0_777 VDD VSS sg13g2_decap_8
XFILLER_75_567 VDD VSS sg13g2_decap_8
XFILLER_90_504 VDD VSS sg13g2_decap_8
XFILLER_29_973 VDD VSS sg13g2_decap_8
X_2196__148 VDD VSS _2196_/RESET_B sg13g2_tiehi
XFILLER_62_206 VDD VSS sg13g2_fill_2
XFILLER_44_921 VDD VSS sg13g2_decap_8
XFILLER_56_770 VDD VSS sg13g2_decap_8
XFILLER_16_623 VDD VSS sg13g2_decap_8
XFILLER_46_63 VDD VSS sg13g2_decap_8
XFILLER_28_483 VDD VSS sg13g2_decap_8
XFILLER_55_280 VDD VSS sg13g2_decap_8
XFILLER_15_133 VDD VSS sg13g2_decap_8
XIO_CORNER_SOUTH_WEST_INST IOVDD IOVSS VDD VSS sg13g2_Corner
XFILLER_43_420 VDD VSS sg13g2_decap_8
XFILLER_71_784 VDD VSS sg13g2_decap_8
XFILLER_102_91 VDD VSS sg13g2_decap_8
XFILLER_44_998 VDD VSS sg13g2_decap_8
XFILLER_31_637 VDD VSS sg13g2_decap_8
XFILLER_12_840 VDD VSS sg13g2_decap_8
XFILLER_50_1017 VDD VSS sg13g2_fill_2
XFILLER_11_350 VDD VSS sg13g2_decap_8
XFILLER_30_147 VDD VSS sg13g2_decap_8
XFILLER_62_84 VDD VSS sg13g2_decap_8
XFILLER_50_1028 VDD VSS sg13g2_fill_1
XFILLER_7_35 VDD VSS sg13g2_decap_8
XFILLER_8_833 VDD VSS sg13g2_decap_8
XFILLER_7_343 VDD VSS sg13g2_decap_8
XFILLER_98_626 VDD VSS sg13g2_decap_8
XFILLER_3_560 VDD VSS sg13g2_decap_8
XFILLER_100_609 VDD VSS sg13g2_decap_8
XFILLER_79_851 VDD VSS sg13g2_fill_2
XFILLER_97_147 VDD VSS sg13g2_decap_4
XFILLER_97_158 VDD VSS sg13g2_fill_1
X_2221_ _2221__98/L_HI VSS VDD _2221_/D _2221_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_87_70 VDD VSS sg13g2_decap_8
XFILLER_79_895 VDD VSS sg13g2_decap_8
XFILLER_112_469 VDD VSS sg13g2_decap_8
XFILLER_66_512 VDD VSS sg13g2_decap_8
XFILLER_38_203 VDD VSS sg13g2_decap_8
X_2152_ _2162_/B _2040_/A _2331_/D VDD VSS sg13g2_nor2b_1
XFILLER_39_759 VDD VSS sg13g2_decap_8
X_2083_ _2083_/A _2089_/S _2083_/Y VDD VSS sg13g2_nor2b_1
XFILLER_93_397 VDD VSS sg13g2_decap_8
XFILLER_35_910 VDD VSS sg13g2_decap_8
XFILLER_19_483 VDD VSS sg13g2_decap_8
XFILLER_81_559 VDD VSS sg13g2_decap_8
XFILLER_62_740 VDD VSS sg13g2_decap_8
XFILLER_34_420 VDD VSS sg13g2_decap_8
XFILLER_46_291 VDD VSS sg13g2_fill_1
XFILLER_35_987 VDD VSS sg13g2_decap_8
XFILLER_99_0 VDD VSS sg13g2_decap_8
XFILLER_50_946 VDD VSS sg13g2_decap_8
XFILLER_22_637 VDD VSS sg13g2_decap_8
XFILLER_61_294 VDD VSS sg13g2_decap_8
XFILLER_34_497 VDD VSS sg13g2_decap_8
XFILLER_21_147 VDD VSS sg13g2_decap_8
X_1936_ VSS VDD _2048_/A _1935_/Y _1936_/Y _1907_/A sg13g2_a21oi_1
XFILLER_107_208 VDD VSS sg13g2_decap_8
XFILLER_107_219 VDD VSS sg13g2_decap_8
X_1867_ _1892_/A _1892_/B _1880_/B _1870_/A VDD VSS sg13g2_nor3_1
X_1798_ _2225_/Q _2217_/Q _1823_/A VDD VSS sg13g2_xor2_1
XFILLER_104_915 VDD VSS sg13g2_decap_8
XFILLER_107_14 VDD VSS sg13g2_decap_8
XFILLER_66_1035 VDD VSS sg13g2_decap_8
XFILLER_27_1008 VDD VSS sg13g2_decap_8
XFILLER_89_659 VDD VSS sg13g2_fill_1
XFILLER_103_458 VDD VSS sg13g2_decap_8
XFILLER_88_147 VDD VSS sg13g2_decap_8
XFILLER_85_810 VDD VSS sg13g2_decap_8
XFILLER_69_372 VDD VSS sg13g2_decap_8
XFILLER_29_203 VDD VSS sg13g2_decap_8
XFILLER_85_887 VDD VSS sg13g2_decap_4
XFILLER_72_504 VDD VSS sg13g2_decap_8
XFILLER_57_567 VDD VSS sg13g2_decap_8
XFILLER_72_515 VDD VSS sg13g2_decap_8
XFILLER_83_28 VDD VSS sg13g2_decap_8
XFILLER_26_910 VDD VSS sg13g2_decap_8
XFILLER_72_559 VDD VSS sg13g2_fill_1
XFILLER_25_420 VDD VSS sg13g2_decap_8
XFILLER_37_280 VDD VSS sg13g2_decap_8
XFILLER_26_987 VDD VSS sg13g2_decap_8
XFILLER_41_902 VDD VSS sg13g2_decap_8
XFILLER_16_77 VDD VSS sg13g2_decap_8
XFILLER_52_261 VDD VSS sg13g2_fill_2
XFILLER_52_250 VDD VSS sg13g2_decap_8
XFILLER_13_637 VDD VSS sg13g2_decap_8
XFILLER_25_497 VDD VSS sg13g2_decap_8
XFILLER_40_412 VDD VSS sg13g2_decap_8
XFILLER_52_283 VDD VSS sg13g2_fill_1
XFILLER_41_979 VDD VSS sg13g2_decap_8
XFILLER_12_147 VDD VSS sg13g2_decap_8
XFILLER_32_21 VDD VSS sg13g2_decap_8
XFILLER_32_98 VDD VSS sg13g2_decap_8
XFILLER_5_847 VDD VSS sg13g2_decap_8
XFILLER_10_1001 VDD VSS sg13g2_decap_8
XFILLER_4_357 VDD VSS sg13g2_decap_8
XFILLER_107_786 VDD VSS sg13g2_decap_8
XFILLER_106_252 VDD VSS sg13g2_decap_8
XFILLER_110_907 VDD VSS sg13g2_decap_8
XFILLER_79_147 VDD VSS sg13g2_decap_8
XFILLER_79_169 VDD VSS sg13g2_decap_8
XFILLER_0_574 VDD VSS sg13g2_decap_8
XFILLER_102_491 VDD VSS sg13g2_decap_8
XFILLER_75_320 VDD VSS sg13g2_decap_8
XFILLER_76_865 VDD VSS sg13g2_decap_8
XFILLER_36_707 VDD VSS sg13g2_decap_8
XFILLER_57_95 VDD VSS sg13g2_decap_4
XFILLER_90_312 VDD VSS sg13g2_decap_8
XFILLER_48_589 VDD VSS sg13g2_decap_8
XFILLER_29_770 VDD VSS sg13g2_decap_8
XFILLER_17_910 VDD VSS sg13g2_decap_8
XFILLER_35_217 VDD VSS sg13g2_decap_8
XFILLER_91_857 VDD VSS sg13g2_decap_8
XFILLER_63_559 VDD VSS sg13g2_decap_8
XFILLER_16_420 VDD VSS sg13g2_decap_8
XFILLER_28_280 VDD VSS sg13g2_decap_8
XFILLER_32_924 VDD VSS sg13g2_decap_8
XFILLER_17_987 VDD VSS sg13g2_decap_8
XFILLER_50_209 VDD VSS sg13g2_decap_8
XFILLER_92_7 VDD VSS sg13g2_decap_8
XFILLER_44_795 VDD VSS sg13g2_decap_4
XFILLER_16_497 VDD VSS sg13g2_decap_8
XFILLER_31_434 VDD VSS sg13g2_decap_8
XFILLER_43_272 VDD VSS sg13g2_decap_8
XFILLER_8_630 VDD VSS sg13g2_decap_8
XFILLER_89_1024 VDD VSS sg13g2_fill_1
X_1721_ _1720_/Y VDD _1721_/Y VSS _1720_/A hold472/X sg13g2_o21ai_1
XFILLER_7_140 VDD VSS sg13g2_decap_8
XFILLER_89_1057 VDD VSS sg13g2_decap_4
X_1652_ _1671_/C _1652_/B _2300_/D VDD VSS sg13g2_nor2_1
X_1583_ _1583_/A _1583_/B _2282_/D VDD VSS sg13g2_nor2_1
XFILLER_99_979 VDD VSS sg13g2_decap_8
XFILLER_101_907 VDD VSS sg13g2_decap_8
XFILLER_98_91 VDD VSS sg13g2_decap_8
XFILLER_86_607 VDD VSS sg13g2_decap_4
XFILLER_112_266 VDD VSS sg13g2_decap_8
XFILLER_58_309 VDD VSS sg13g2_decap_8
XFILLER_79_692 VDD VSS sg13g2_decap_8
XFILLER_100_439 VDD VSS sg13g2_decap_4
X_2204_ _2204_/RESET_B VSS VDD _2204_/D _2204_/Q clkload4/A sg13g2_dfrbpq_1
X_2135_ _2135_/A _2135_/B _2370_/D VDD VSS sg13g2_nor2_1
XFILLER_94_662 VDD VSS sg13g2_decap_8
XFILLER_94_640 VDD VSS sg13g2_fill_1
XFILLER_82_813 VDD VSS sg13g2_decap_8
XFILLER_39_556 VDD VSS sg13g2_decap_8
XFILLER_27_707 VDD VSS sg13g2_decap_8
XFILLER_14_0 VDD VSS sg13g2_decap_8
XFILLER_96_1039 VDD VSS sg13g2_decap_8
XFILLER_81_312 VDD VSS sg13g2_decap_8
XFILLER_93_161 VDD VSS sg13g2_decap_4
XFILLER_26_217 VDD VSS sg13g2_decap_8
XFILLER_82_879 VDD VSS sg13g2_decap_8
X_2066_ _2338_/D _2066_/A _2066_/B VDD VSS sg13g2_nand2_1
XFILLER_19_280 VDD VSS sg13g2_decap_8
XFILLER_23_924 VDD VSS sg13g2_decap_8
XFILLER_35_784 VDD VSS sg13g2_decap_8
XFILLER_41_209 VDD VSS sg13g2_decap_8
XFILLER_22_434 VDD VSS sg13g2_decap_8
XFILLER_34_294 VDD VSS sg13g2_decap_8
XFILLER_33_1001 VDD VSS sg13g2_decap_8
XFILLER_50_798 VDD VSS sg13g2_decap_8
X_1919_ _1919_/B _1919_/A _1924_/A VDD VSS sg13g2_xor2_1
XFILLER_108_528 VDD VSS sg13g2_decap_8
XFILLER_89_412 VDD VSS sg13g2_decap_8
XFILLER_78_28 VDD VSS sg13g2_decap_8
XFILLER_104_778 VDD VSS sg13g2_decap_8
XFILLER_77_607 VDD VSS sg13g2_decap_8
XFILLER_49_309 VDD VSS sg13g2_decap_8
XFILLER_98_990 VDD VSS sg13g2_decap_8
XFILLER_103_277 VDD VSS sg13g2_decap_8
XFILLER_40_1005 VDD VSS sg13g2_decap_8
XFILLER_100_973 VDD VSS sg13g2_decap_8
XFILLER_94_49 VDD VSS sg13g2_decap_8
XFILLER_18_707 VDD VSS sg13g2_decap_8
XFILLER_73_846 VDD VSS sg13g2_decap_8
XFILLER_72_301 VDD VSS sg13g2_decap_8
XFILLER_72_312 VDD VSS sg13g2_fill_1
XFILLER_17_217 VDD VSS sg13g2_decap_8
XFILLER_27_21 VDD VSS sg13g2_decap_8
XFILLER_45_504 VDD VSS sg13g2_decap_8
XFILLER_72_345 VDD VSS sg13g2_decap_8
XFILLER_57_397 VDD VSS sg13g2_decap_8
XFILLER_26_784 VDD VSS sg13g2_decap_8
XFILLER_14_924 VDD VSS sg13g2_decap_8
XFILLER_27_98 VDD VSS sg13g2_decap_8
XFILLER_13_434 VDD VSS sg13g2_decap_8
XFILLER_25_294 VDD VSS sg13g2_decap_8
XFILLER_41_776 VDD VSS sg13g2_decap_8
XFILLER_43_42 VDD VSS sg13g2_decap_8
XFILLER_9_427 VDD VSS sg13g2_decap_8
XFILLER_40_286 VDD VSS sg13g2_fill_1
X_2226__88 VDD VSS _2226__88/L_HI sg13g2_tiehi
XFILLER_99_209 VDD VSS sg13g2_fill_1
XFILLER_5_644 VDD VSS sg13g2_decap_8
XFILLER_107_583 VDD VSS sg13g2_decap_8
XFILLER_4_14 VDD VSS sg13g2_decap_8
XFILLER_4_154 VDD VSS sg13g2_decap_8
XFILLER_96_927 VDD VSS sg13g2_fill_2
XFILLER_110_704 VDD VSS sg13g2_decap_8
XFILLER_68_629 VDD VSS sg13g2_decap_4
XFILLER_1_861 VDD VSS sg13g2_decap_8
XFILLER_95_448 VDD VSS sg13g2_decap_8
XFILLER_49_843 VDD VSS sg13g2_fill_1
XFILLER_49_832 VDD VSS sg13g2_decap_8
XFILLER_0_371 VDD VSS sg13g2_decap_8
XFILLER_64_802 VDD VSS sg13g2_decap_8
XFILLER_49_876 VDD VSS sg13g2_decap_8
XFILLER_75_161 VDD VSS sg13g2_decap_4
XFILLER_36_504 VDD VSS sg13g2_decap_8
XFILLER_63_345 VDD VSS sg13g2_decap_8
XFILLER_1_1043 VDD VSS sg13g2_decap_8
XFILLER_95_1050 VDD VSS sg13g2_decap_8
XFILLER_91_676 VDD VSS sg13g2_decap_8
XFILLER_90_153 VDD VSS sg13g2_decap_8
XFILLER_56_1012 VDD VSS sg13g2_fill_1
XFILLER_44_592 VDD VSS sg13g2_decap_8
XFILLER_32_721 VDD VSS sg13g2_decap_8
XFILLER_17_784 VDD VSS sg13g2_decap_8
XFILLER_16_294 VDD VSS sg13g2_decap_8
XFILLER_17_1029 VDD VSS sg13g2_decap_8
XFILLER_31_231 VDD VSS sg13g2_decap_8
XFILLER_32_798 VDD VSS sg13g2_decap_8
XFILLER_20_938 VDD VSS sg13g2_decap_8
X_1704_ _1705_/B _1704_/A _1709_/A VDD VSS sg13g2_xnor2_1
XFILLER_9_994 VDD VSS sg13g2_decap_8
X_1635_ _1634_/Y VDD _1635_/Y VSS _1634_/A hold542/X sg13g2_o21ai_1
X_1566_ _1565_/Y VDD _1566_/Y VSS _1573_/A1 hold421/X sg13g2_o21ai_1
XFILLER_99_787 VDD VSS sg13g2_decap_8
XFILLER_98_253 VDD VSS sg13g2_decap_8
XFILLER_101_726 VDD VSS sg13g2_decap_8
XFILLER_86_426 VDD VSS sg13g2_decap_8
XFILLER_58_128 VDD VSS sg13g2_decap_8
X_1497_ _1497_/A _1497_/B _1497_/C _1497_/Y VDD VSS sg13g2_nor3_1
XFILLER_100_247 VDD VSS sg13g2_decap_8
XFILLER_39_331 VDD VSS sg13g2_decap_8
XFILLER_67_684 VDD VSS sg13g2_decap_8
XFILLER_27_504 VDD VSS sg13g2_decap_8
XFILLER_82_632 VDD VSS sg13g2_decap_8
X_2118_ hold530/X VDD _2118_/Y VSS _2144_/S0 hold394/X sg13g2_o21ai_1
XFILLER_55_846 VDD VSS sg13g2_decap_8
XFILLER_54_334 VDD VSS sg13g2_decap_8
X_2049_ _1936_/Y _1908_/A _2069_/S _2049_/X VDD VSS sg13g2_mux2_1
XFILLER_81_164 VDD VSS sg13g2_decap_8
Xfanout13 _2007_/B _2071_/B VDD VSS sg13g2_buf_1
XFILLER_81_197 VDD VSS sg13g2_fill_2
XFILLER_81_175 VDD VSS sg13g2_fill_2
XFILLER_35_581 VDD VSS sg13g2_decap_8
XFILLER_23_721 VDD VSS sg13g2_decap_8
Xfanout35 fanout40/X _1342_/A2 VDD VSS sg13g2_buf_1
Xfanout46 _2311_/Q _1677_/A VDD VSS sg13g2_buf_1
Xfanout24 _1465_/Y _1481_/A2 VDD VSS sg13g2_buf_1
XFILLER_22_231 VDD VSS sg13g2_decap_8
Xfanout68 _1228_/A _1671_/C VDD VSS sg13g2_buf_1
XFILLER_23_798 VDD VSS sg13g2_decap_8
XFILLER_11_938 VDD VSS sg13g2_decap_8
Xfanout57 _1634_/A _1638_/S VDD VSS sg13g2_buf_1
XFILLER_10_448 VDD VSS sg13g2_decap_8
XFILLER_13_56 VDD VSS sg13g2_decap_8
XFILLER_109_826 VDD VSS sg13g2_decap_8
XFILLER_108_347 VDD VSS sg13g2_decap_8
XFILLER_89_49 VDD VSS sg13g2_decap_8
Xhold471 _2224_/Q VDD VSS hold471/X sg13g2_dlygate4sd3_1
XFILLER_104_531 VDD VSS sg13g2_decap_8
Xhold460 _2251_/Q VDD VSS _1463_/A sg13g2_dlygate4sd3_1
XFILLER_2_658 VDD VSS sg13g2_decap_8
XFILLER_78_916 VDD VSS sg13g2_decap_8
Xhold493 _2233_/Q VDD VSS _1424_/A sg13g2_dlygate4sd3_1
Xhold482 _2248_/Q VDD VSS _1457_/A sg13g2_dlygate4sd3_1
XFILLER_89_286 VDD VSS sg13g2_decap_8
XFILLER_77_426 VDD VSS sg13g2_decap_4
XFILLER_1_168 VDD VSS sg13g2_decap_8
XFILLER_93_908 VDD VSS sg13g2_fill_2
XFILLER_58_651 VDD VSS sg13g2_decap_8
XFILLER_38_42 VDD VSS sg13g2_decap_8
XFILLER_79_1001 VDD VSS sg13g2_decap_8
XFILLER_46_824 VDD VSS sg13g2_decap_8
XFILLER_18_504 VDD VSS sg13g2_decap_8
XFILLER_57_150 VDD VSS sg13g2_decap_8
XFILLER_45_301 VDD VSS sg13g2_decap_8
XFILLER_57_172 VDD VSS sg13g2_decap_8
XFILLER_33_518 VDD VSS sg13g2_decap_8
XFILLER_72_175 VDD VSS sg13g2_decap_8
XFILLER_26_581 VDD VSS sg13g2_decap_8
XFILLER_14_721 VDD VSS sg13g2_decap_8
XFILLER_60_359 VDD VSS sg13g2_decap_8
XFILLER_13_231 VDD VSS sg13g2_decap_8
XFILLER_54_85 VDD VSS sg13g2_decap_8
XFILLER_9_224 VDD VSS sg13g2_decap_8
XFILLER_14_798 VDD VSS sg13g2_decap_8
XFILLER_110_91 VDD VSS sg13g2_decap_8
XFILLER_103_1043 VDD VSS sg13g2_decap_8
XFILLER_70_84 VDD VSS sg13g2_decap_8
XFILLER_6_931 VDD VSS sg13g2_decap_8
XFILLER_86_1005 VDD VSS sg13g2_fill_1
XFILLER_5_441 VDD VSS sg13g2_decap_8
XFILLER_55_7 VDD VSS sg13g2_decap_8
XFILLER_108_892 VDD VSS sg13g2_decap_8
X_1420_ _1420_/Y _1420_/A _1426_/B VDD VSS sg13g2_nand2_1
X_1351_ VDD _2204_/D _1351_/A VSS sg13g2_inv_1
XFILLER_96_735 VDD VSS sg13g2_decap_8
XFILLER_110_501 VDD VSS sg13g2_decap_8
XFILLER_96_768 VDD VSS sg13g2_decap_8
XFILLER_95_234 VDD VSS sg13g2_decap_8
XFILLER_23_1022 VDD VSS sg13g2_decap_8
X_1282_ _1282_/Y _1482_/B1 hold318/X _1482_/A2 _2375_/Q VDD VSS sg13g2_a22oi_1
XFILLER_68_448 VDD VSS sg13g2_fill_2
XFILLER_68_459 VDD VSS sg13g2_decap_8
XFILLER_77_993 VDD VSS sg13g2_decap_8
XFILLER_110_578 VDD VSS sg13g2_decap_8
XFILLER_95_70 VDD VSS sg13g2_decap_8
XFILLER_49_662 VDD VSS sg13g2_decap_8
XFILLER_48_161 VDD VSS sg13g2_decap_8
XFILLER_55_109 VDD VSS sg13g2_decap_8
XFILLER_36_301 VDD VSS sg13g2_decap_8
XFILLER_110_1047 VDD VSS sg13g2_decap_8
XFILLER_37_868 VDD VSS sg13g2_decap_8
XFILLER_92_974 VDD VSS sg13g2_fill_2
XFILLER_91_440 VDD VSS sg13g2_decap_8
XFILLER_64_676 VDD VSS sg13g2_decap_8
XFILLER_63_131 VDD VSS sg13g2_decap_8
XFILLER_24_518 VDD VSS sg13g2_decap_8
XFILLER_36_378 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_52_838 VDD VSS sg13g2_decap_8
XFILLER_52_849 VDD VSS sg13g2_decap_8
XFILLER_51_326 VDD VSS sg13g2_decap_8
XFILLER_17_581 VDD VSS sg13g2_decap_8
XFILLER_60_893 VDD VSS sg13g2_decap_8
XFILLER_81_0 VDD VSS sg13g2_decap_8
XFILLER_32_595 VDD VSS sg13g2_decap_8
XFILLER_20_735 VDD VSS sg13g2_decap_8
XFILLER_30_1015 VDD VSS sg13g2_decap_8
XFILLER_9_791 VDD VSS sg13g2_decap_8
XFILLER_106_818 VDD VSS sg13g2_decap_8
X_1618_ _1619_/B _1618_/A _1623_/A VDD VSS sg13g2_xnor2_1
XFILLER_99_562 VDD VSS sg13g2_decap_8
XFILLER_59_404 VDD VSS sg13g2_decap_8
XFILLER_87_724 VDD VSS sg13g2_decap_8
X_1549_ _1556_/S0 _2238_/Q _2230_/Q _2222_/Q _2214_/Q _1589_/B _1550_/A VDD VSS sg13g2_mux4_1
XFILLER_86_223 VDD VSS sg13g2_decap_8
XFILLER_59_426 VDD VSS sg13g2_decap_8
XFILLER_101_534 VDD VSS sg13g2_decap_8
XFILLER_39_161 VDD VSS sg13g2_decap_8
XFILLER_27_301 VDD VSS sg13g2_decap_8
XFILLER_28_868 VDD VSS sg13g2_decap_8
XFILLER_54_120 VDD VSS sg13g2_decap_8
XFILLER_83_974 VDD VSS sg13g2_decap_8
XFILLER_15_518 VDD VSS sg13g2_decap_8
XFILLER_27_378 VDD VSS sg13g2_decap_8
XFILLER_91_28 VDD VSS sg13g2_decap_8
XFILLER_43_849 VDD VSS sg13g2_decap_8
XFILLER_54_175 VDD VSS sg13g2_decap_8
XFILLER_70_668 VDD VSS sg13g2_decap_8
XFILLER_23_595 VDD VSS sg13g2_decap_8
XFILLER_11_735 VDD VSS sg13g2_decap_8
XFILLER_24_77 VDD VSS sg13g2_decap_8
XFILLER_50_381 VDD VSS sg13g2_decap_8
XFILLER_109_623 VDD VSS sg13g2_decap_8
XFILLER_10_245 VDD VSS sg13g2_decap_8
XFILLER_7_728 VDD VSS sg13g2_decap_8
XFILLER_108_133 VDD VSS sg13g2_decap_8
XFILLER_6_238 VDD VSS sg13g2_decap_8
XFILLER_40_21 VDD VSS sg13g2_decap_8
XFILLER_105_840 VDD VSS sg13g2_decap_8
XFILLER_3_945 VDD VSS sg13g2_decap_8
XFILLER_40_98 VDD VSS sg13g2_decap_8
XFILLER_2_455 VDD VSS sg13g2_decap_8
X_2242__258 VDD VSS _2242_/RESET_B sg13g2_tiehi
XFILLER_49_63 VDD VSS sg13g2_decap_8
XFILLER_78_768 VDD VSS sg13g2_decap_8
XFILLER_77_256 VDD VSS sg13g2_decap_4
XFILLER_49_74 VDD VSS sg13g2_fill_1
XFILLER_49_96 VDD VSS sg13g2_decap_8
XFILLER_93_738 VDD VSS sg13g2_decap_8
XFILLER_59_971 VDD VSS sg13g2_decap_8
XFILLER_18_301 VDD VSS sg13g2_decap_8
XFILLER_105_91 VDD VSS sg13g2_decap_8
XFILLER_46_621 VDD VSS sg13g2_decap_8
XFILLER_34_805 VDD VSS sg13g2_decap_8
XFILLER_19_868 VDD VSS sg13g2_decap_8
XFILLER_65_73 VDD VSS sg13g2_decap_8
XFILLER_73_484 VDD VSS sg13g2_decap_8
XFILLER_18_378 VDD VSS sg13g2_decap_8
XFILLER_33_315 VDD VSS sg13g2_decap_8
XFILLER_45_175 VDD VSS sg13g2_decap_8
XFILLER_92_1031 VDD VSS sg13g2_decap_8
X_2175__190 VDD VSS _2175_/RESET_B sg13g2_tiehi
XFILLER_53_1004 VDD VSS sg13g2_decap_8
XFILLER_42_882 VDD VSS sg13g2_decap_8
XFILLER_14_595 VDD VSS sg13g2_decap_8
XFILLER_41_381 VDD VSS sg13g2_decap_8
XFILLER_69_713 VDD VSS sg13g2_decap_8
X_1403_ _1404_/A _1392_/Y hold471/X _1392_/B _1382_/A VDD VSS sg13g2_a22oi_1
XFILLER_96_521 VDD VSS sg13g2_decap_8
XFILLER_111_854 VDD VSS sg13g2_decap_8
X_1334_ _1334_/Y _1342_/B1 hold401/X _1342_/A2 _2330_/Q VDD VSS sg13g2_a22oi_1
XFILLER_57_908 VDD VSS sg13g2_decap_8
XFILLER_110_375 VDD VSS sg13g2_decap_8
X_1265_ _2150_/A _1265_/B _1265_/X VDD VSS sg13g2_and2_1
XFILLER_65_930 VDD VSS sg13g2_decap_8
XFILLER_37_665 VDD VSS sg13g2_decap_8
XFILLER_25_805 VDD VSS sg13g2_decap_8
XFILLER_64_451 VDD VSS sg13g2_decap_8
X_1196_ VDD _1196_/Y _1196_/A VSS sg13g2_inv_1
XFILLER_52_624 VDD VSS sg13g2_decap_8
XFILLER_51_112 VDD VSS sg13g2_decap_8
XFILLER_24_315 VDD VSS sg13g2_decap_8
XFILLER_36_175 VDD VSS sg13g2_decap_8
XFILLER_80_966 VDD VSS sg13g2_decap_8
XFILLER_101_49 VDD VSS sg13g2_decap_8
XFILLER_33_882 VDD VSS sg13g2_decap_8
XFILLER_20_532 VDD VSS sg13g2_decap_8
XFILLER_32_392 VDD VSS sg13g2_decap_8
XFILLER_106_615 VDD VSS sg13g2_decap_8
XFILLER_10_35 VDD VSS sg13g2_decap_8
XFILLER_105_147 VDD VSS sg13g2_fill_2
XFILLER_102_832 VDD VSS sg13g2_decap_8
XFILLER_87_521 VDD VSS sg13g2_decap_4
XFILLER_86_28 VDD VSS sg13g2_decap_8
XFILLER_59_201 VDD VSS sg13g2_decap_8
XFILLER_87_532 VDD VSS sg13g2_fill_1
XFILLER_48_908 VDD VSS sg13g2_decap_8
XFILLER_0_959 VDD VSS sg13g2_decap_8
XFILLER_87_576 VDD VSS sg13g2_decap_8
XFILLER_75_749 VDD VSS sg13g2_decap_8
XFILLER_101_386 VDD VSS sg13g2_decap_8
XFILLER_74_237 VDD VSS sg13g2_decap_8
XFILLER_56_941 VDD VSS sg13g2_decap_8
XFILLER_19_77 VDD VSS sg13g2_decap_8
XFILLER_71_900 VDD VSS sg13g2_decap_8
XFILLER_28_665 VDD VSS sg13g2_decap_8
XFILLER_16_805 VDD VSS sg13g2_decap_8
XFILLER_70_421 VDD VSS sg13g2_fill_1
XFILLER_55_473 VDD VSS sg13g2_decap_8
XFILLER_15_315 VDD VSS sg13g2_decap_8
XFILLER_35_21 VDD VSS sg13g2_decap_8
XFILLER_42_112 VDD VSS sg13g2_decap_8
XFILLER_27_175 VDD VSS sg13g2_decap_8
XFILLER_71_977 VDD VSS sg13g2_decap_8
XFILLER_82_292 VDD VSS sg13g2_decap_8
XFILLER_43_646 VDD VSS sg13g2_decap_8
XIO_BOND_in_valid_pad in_valid_PAD bondpad_70x70
XFILLER_31_819 VDD VSS sg13g2_decap_8
XFILLER_24_882 VDD VSS sg13g2_decap_8
XFILLER_35_98 VDD VSS sg13g2_decap_8
XFILLER_42_156 VDD VSS sg13g2_decap_8
XFILLER_70_498 VDD VSS sg13g2_decap_8
XFILLER_11_532 VDD VSS sg13g2_decap_8
XFILLER_23_392 VDD VSS sg13g2_decap_8
XFILLER_30_329 VDD VSS sg13g2_decap_8
XFILLER_109_420 VDD VSS sg13g2_decap_8
XFILLER_7_525 VDD VSS sg13g2_decap_8
XFILLER_13_1043 VDD VSS sg13g2_decap_8
XFILLER_109_497 VDD VSS sg13g2_decap_8
XFILLER_83_1008 VDD VSS sg13g2_decap_4
XFILLER_3_742 VDD VSS sg13g2_decap_8
XFILLER_97_329 VDD VSS sg13g2_decap_8
XFILLER_2_252 VDD VSS sg13g2_decap_8
XFILLER_38_418 VDD VSS sg13g2_decap_8
XFILLER_65_226 VDD VSS sg13g2_decap_8
XFILLER_18_7 VDD VSS sg13g2_decap_8
XFILLER_93_579 VDD VSS sg13g2_decap_8
XFILLER_81_708 VDD VSS sg13g2_decap_8
XFILLER_47_985 VDD VSS sg13g2_decap_8
XFILLER_19_665 VDD VSS sg13g2_decap_8
XFILLER_20_1036 VDD VSS sg13g2_decap_8
XFILLER_74_793 VDD VSS sg13g2_decap_8
XFILLER_73_270 VDD VSS sg13g2_decap_8
XFILLER_34_602 VDD VSS sg13g2_decap_8
XFILLER_18_175 VDD VSS sg13g2_decap_8
XFILLER_73_292 VDD VSS sg13g2_decap_8
XFILLER_73_281 VDD VSS sg13g2_fill_2
XFILLER_61_432 VDD VSS sg13g2_decap_8
XFILLER_33_112 VDD VSS sg13g2_decap_8
XFILLER_62_999 VDD VSS sg13g2_decap_8
XFILLER_34_679 VDD VSS sg13g2_decap_8
XFILLER_22_819 VDD VSS sg13g2_decap_8
XFILLER_15_882 VDD VSS sg13g2_decap_8
X_1952_ _1952_/B _1952_/A _1953_/A VDD VSS sg13g2_xor2_1
XFILLER_61_498 VDD VSS sg13g2_decap_8
XFILLER_14_392 VDD VSS sg13g2_decap_8
XFILLER_21_329 VDD VSS sg13g2_decap_8
XFILLER_33_189 VDD VSS sg13g2_decap_8
X_1883_ _1879_/B _1879_/A _1882_/Y _1972_/A VDD VSS sg13g2_a21o_1
XFILLER_30_896 VDD VSS sg13g2_decap_8
XFILLER_44_0 VDD VSS sg13g2_decap_8
XFILLER_29_1050 VDD VSS sg13g2_decap_8
XFILLER_111_651 VDD VSS sg13g2_decap_8
XFILLER_97_874 VDD VSS sg13g2_decap_8
XFILLER_69_565 VDD VSS sg13g2_decap_8
X_2366_ _2366_/RESET_B VSS VDD _2366_/D _2366_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_57_716 VDD VSS sg13g2_decap_8
XFILLER_5_1008 VDD VSS sg13g2_decap_8
XFILLER_110_161 VDD VSS sg13g2_decap_8
X_1317_ VDD _2188_/D _1317_/A VSS sg13g2_inv_1
X_2297_ _2297_/RESET_B VSS VDD _2297_/D _2297_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_2_91 VDD VSS sg13g2_decap_8
X_1248_ _1248_/B _1248_/C _1248_/A _1249_/C VDD VSS sg13g2_nand3_1
XFILLER_71_229 VDD VSS sg13g2_decap_8
XFILLER_53_933 VDD VSS sg13g2_decap_4
XFILLER_38_996 VDD VSS sg13g2_decap_8
XFILLER_53_911 VDD VSS sg13g2_decap_8
XFILLER_25_602 VDD VSS sg13g2_decap_8
XFILLER_52_410 VDD VSS sg13g2_decap_8
XFILLER_37_462 VDD VSS sg13g2_decap_8
XFILLER_53_955 VDD VSS sg13g2_decap_8
XFILLER_53_944 VDD VSS sg13g2_fill_2
XFILLER_24_112 VDD VSS sg13g2_decap_8
XFILLER_80_774 VDD VSS sg13g2_decap_8
XFILLER_40_627 VDD VSS sg13g2_decap_8
XFILLER_25_679 VDD VSS sg13g2_decap_8
XFILLER_13_819 VDD VSS sg13g2_decap_8
XFILLER_36_1043 VDD VSS sg13g2_decap_8
XFILLER_12_329 VDD VSS sg13g2_decap_8
XFILLER_24_189 VDD VSS sg13g2_decap_8
XFILLER_21_896 VDD VSS sg13g2_decap_8
XFILLER_4_539 VDD VSS sg13g2_decap_8
XFILLER_21_56 VDD VSS sg13g2_decap_8
XFILLER_107_968 VDD VSS sg13g2_decap_8
XFILLER_106_456 VDD VSS sg13g2_decap_8
XIO_BOND_in_data_pads\[2\].in_data_pad in_data_PADs[2] bondpad_70x70
XFILLER_97_49 VDD VSS sg13g2_decap_8
XFILLER_88_830 VDD VSS sg13g2_decap_8
XFILLER_43_1003 VDD VSS sg13g2_decap_8
XFILLER_0_756 VDD VSS sg13g2_decap_8
XFILLER_102_673 VDD VSS sg13g2_decap_4
XFILLER_102_684 VDD VSS sg13g2_decap_4
XFILLER_101_183 VDD VSS sg13g2_fill_2
XFILLER_87_395 VDD VSS sg13g2_decap_8
XFILLER_75_535 VDD VSS sg13g2_decap_8
XFILLER_29_952 VDD VSS sg13g2_decap_8
XFILLER_44_900 VDD VSS sg13g2_decap_8
XFILLER_46_42 VDD VSS sg13g2_decap_8
XFILLER_62_218 VDD VSS sg13g2_fill_1
XFILLER_16_602 VDD VSS sg13g2_decap_8
XFILLER_28_462 VDD VSS sg13g2_decap_8
XFILLER_90_549 VDD VSS sg13g2_decap_8
XFILLER_71_741 VDD VSS sg13g2_decap_8
XFILLER_44_977 VDD VSS sg13g2_decap_8
XFILLER_15_112 VDD VSS sg13g2_decap_8
XFILLER_71_763 VDD VSS sg13g2_decap_8
XFILLER_70_262 VDD VSS sg13g2_fill_1
XFILLER_102_70 VDD VSS sg13g2_decap_8
XFILLER_31_616 VDD VSS sg13g2_decap_8
XFILLER_16_679 VDD VSS sg13g2_decap_8
XFILLER_15_189 VDD VSS sg13g2_decap_8
XFILLER_30_126 VDD VSS sg13g2_decap_8
XFILLER_62_63 VDD VSS sg13g2_decap_8
XFILLER_43_498 VDD VSS sg13g2_fill_1
XFILLER_8_812 VDD VSS sg13g2_decap_8
XFILLER_7_322 VDD VSS sg13g2_decap_8
XFILLER_7_14 VDD VSS sg13g2_decap_8
XFILLER_12_896 VDD VSS sg13g2_decap_8
XFILLER_8_889 VDD VSS sg13g2_decap_8
XFILLER_109_261 VDD VSS sg13g2_fill_2
XFILLER_109_272 VDD VSS sg13g2_decap_8
XFILLER_7_399 VDD VSS sg13g2_decap_8
XFILLER_112_448 VDD VSS sg13g2_decap_8
XFILLER_97_126 VDD VSS sg13g2_decap_8
X_2220_ _2220_/RESET_B VSS VDD _2220_/D _2220_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_94_822 VDD VSS sg13g2_decap_8
X_2151_ _2156_/A _2040_/A _2330_/D VDD VSS sg13g2_nor2b_1
XFILLER_93_310 VDD VSS sg13g2_decap_8
XFILLER_39_738 VDD VSS sg13g2_decap_8
X_2082_ _2082_/Y _2082_/B _2081_/Y VDD VSS sg13g2_nand2b_1
XFILLER_66_568 VDD VSS sg13g2_decap_8
XFILLER_54_719 VDD VSS sg13g2_decap_4
XFILLER_38_259 VDD VSS sg13g2_decap_8
XFILLER_94_899 VDD VSS sg13g2_decap_8
XFILLER_93_376 VDD VSS sg13g2_decap_8
XFILLER_81_538 VDD VSS sg13g2_decap_8
XFILLER_47_771 VDD VSS sg13g2_decap_8
XFILLER_47_782 VDD VSS sg13g2_fill_1
XFILLER_19_462 VDD VSS sg13g2_decap_8
XFILLER_35_966 VDD VSS sg13g2_decap_8
XFILLER_46_270 VDD VSS sg13g2_decap_8
XFILLER_50_925 VDD VSS sg13g2_decap_8
XFILLER_22_616 VDD VSS sg13g2_decap_8
XFILLER_34_476 VDD VSS sg13g2_decap_8
XFILLER_61_273 VDD VSS sg13g2_decap_8
XFILLER_21_126 VDD VSS sg13g2_decap_8
X_1935_ VDD _1935_/Y _1935_/A VSS sg13g2_inv_1
XFILLER_30_693 VDD VSS sg13g2_decap_8
X_1866_ _1866_/A _1866_/B _1880_/B VDD VSS sg13g2_and2_1
X_1797_ _1797_/Y _2225_/Q _2217_/Q VDD VSS sg13g2_nand2b_1
XFILLER_66_1014 VDD VSS sg13g2_decap_8
XFILLER_89_638 VDD VSS sg13g2_decap_8
XFILLER_103_404 VDD VSS sg13g2_fill_1
X_2262__228 VDD VSS _2262_/RESET_B sg13g2_tiehi
XFILLER_103_437 VDD VSS sg13g2_decap_8
XFILLER_88_126 VDD VSS sg13g2_decap_8
XFILLER_69_362 VDD VSS sg13g2_decap_4
XFILLER_97_682 VDD VSS sg13g2_fill_2
XFILLER_84_321 VDD VSS sg13g2_decap_4
X_2349_ _2349_/RESET_B VSS VDD _2349_/D _2349_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_57_535 VDD VSS sg13g2_fill_2
XFILLER_85_866 VDD VSS sg13g2_decap_8
XFILLER_45_708 VDD VSS sg13g2_fill_2
XFILLER_29_259 VDD VSS sg13g2_decap_8
XFILLER_38_793 VDD VSS sg13g2_decap_8
XFILLER_44_207 VDD VSS sg13g2_decap_8
XFILLER_26_966 VDD VSS sg13g2_decap_8
XFILLER_53_774 VDD VSS sg13g2_fill_1
XFILLER_16_56 VDD VSS sg13g2_decap_8
XFILLER_13_616 VDD VSS sg13g2_decap_8
XFILLER_25_476 VDD VSS sg13g2_decap_8
XFILLER_41_958 VDD VSS sg13g2_decap_8
XFILLER_12_126 VDD VSS sg13g2_decap_8
XFILLER_9_609 VDD VSS sg13g2_decap_8
XFILLER_40_468 VDD VSS sg13g2_decap_4
XFILLER_8_119 VDD VSS sg13g2_decap_8
XFILLER_21_693 VDD VSS sg13g2_decap_8
XFILLER_32_77 VDD VSS sg13g2_decap_8
XFILLER_5_826 VDD VSS sg13g2_decap_8
XFILLER_107_765 VDD VSS sg13g2_decap_8
XFILLER_106_231 VDD VSS sg13g2_decap_8
XFILLER_4_336 VDD VSS sg13g2_decap_8
XFILLER_10_1057 VDD VSS sg13g2_decap_4
XFILLER_79_126 VDD VSS sg13g2_decap_8
XFILLER_0_553 VDD VSS sg13g2_decap_8
XFILLER_88_693 VDD VSS sg13g2_decap_8
XFILLER_76_844 VDD VSS sg13g2_decap_8
XFILLER_102_470 VDD VSS sg13g2_decap_8
XFILLER_48_568 VDD VSS sg13g2_decap_8
XFILLER_57_74 VDD VSS sg13g2_decap_8
XFILLER_91_847 VDD VSS sg13g2_fill_1
XFILLER_63_538 VDD VSS sg13g2_decap_8
XFILLER_90_357 VDD VSS sg13g2_fill_2
XFILLER_17_966 VDD VSS sg13g2_decap_8
XFILLER_44_774 VDD VSS sg13g2_decap_8
XFILLER_32_903 VDD VSS sg13g2_decap_8
XFILLER_16_476 VDD VSS sg13g2_decap_8
XFILLER_43_251 VDD VSS sg13g2_decap_8
XFILLER_71_571 VDD VSS sg13g2_fill_2
XFILLER_73_84 VDD VSS sg13g2_decap_8
XFILLER_31_413 VDD VSS sg13g2_decap_8
XFILLER_85_7 VDD VSS sg13g2_decap_8
XFILLER_40_991 VDD VSS sg13g2_decap_8
XFILLER_89_1036 VDD VSS sg13g2_decap_8
XFILLER_89_1003 VDD VSS sg13g2_decap_8
X_1720_ _1720_/Y _1720_/A _1720_/B VDD VSS sg13g2_nand2_1
XFILLER_12_693 VDD VSS sg13g2_decap_8
X_1651_ _1651_/Y _1646_/Y _1650_/X hold437/X _1671_/B VDD VSS sg13g2_a22oi_1
XFILLER_8_686 VDD VSS sg13g2_decap_8
XFILLER_7_196 VDD VSS sg13g2_decap_8
XFILLER_98_70 VDD VSS sg13g2_decap_8
X_1582_ _1582_/Y _1527_/Y _1581_/Y hold511/X _1190_/Y VDD VSS sg13g2_a22oi_1
XFILLER_99_958 VDD VSS sg13g2_decap_8
XFILLER_98_446 VDD VSS sg13g2_fill_2
XFILLER_112_245 VDD VSS sg13g2_decap_8
XFILLER_79_671 VDD VSS sg13g2_decap_8
X_2203_ _2203_/RESET_B VSS VDD _2203_/D _2203_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_513 VDD VSS sg13g2_decap_8
X_2134_ _2138_/B1 VDD _2135_/B VSS _2142_/A1 hold535/X sg13g2_o21ai_1
XFILLER_78_192 VDD VSS sg13g2_decap_8
XFILLER_93_140 VDD VSS sg13g2_decap_8
XFILLER_54_516 VDD VSS sg13g2_decap_8
X_2065_ _2071_/B _2065_/C _2071_/A _2066_/B VDD VSS sg13g2_nand3_1
XFILLER_81_368 VDD VSS sg13g2_fill_2
XFILLER_35_763 VDD VSS sg13g2_decap_8
XFILLER_23_903 VDD VSS sg13g2_decap_8
XFILLER_50_711 VDD VSS sg13g2_decap_8
XFILLER_22_413 VDD VSS sg13g2_decap_8
XFILLER_34_273 VDD VSS sg13g2_decap_8
XFILLER_50_777 VDD VSS sg13g2_decap_8
XFILLER_31_980 VDD VSS sg13g2_decap_8
X_1918_ _1919_/A _1919_/B _1918_/X VDD VSS sg13g2_and2_1
XFILLER_33_1057 VDD VSS sg13g2_decap_4
XFILLER_30_490 VDD VSS sg13g2_decap_8
X_1849_ VSS VDD _1846_/Y _1848_/A _1863_/A _1850_/B sg13g2_a21oi_1
XFILLER_104_757 VDD VSS sg13g2_decap_8
XFILLER_103_256 VDD VSS sg13g2_decap_8
XFILLER_69_170 VDD VSS sg13g2_decap_8
XFILLER_100_952 VDD VSS sg13g2_decap_8
XFILLER_73_803 VDD VSS sg13g2_fill_2
XFILLER_94_28 VDD VSS sg13g2_decap_8
XFILLER_85_696 VDD VSS sg13g2_decap_8
XFILLER_84_184 VDD VSS sg13g2_decap_8
XFILLER_38_590 VDD VSS sg13g2_decap_8
XFILLER_27_77 VDD VSS sg13g2_decap_8
XFILLER_26_763 VDD VSS sg13g2_decap_8
XFILLER_14_903 VDD VSS sg13g2_decap_8
XFILLER_13_413 VDD VSS sg13g2_decap_8
XFILLER_43_21 VDD VSS sg13g2_decap_8
XFILLER_25_273 VDD VSS sg13g2_decap_8
XFILLER_40_210 VDD VSS sg13g2_decap_8
XFILLER_80_390 VDD VSS sg13g2_decap_8
XFILLER_41_755 VDD VSS sg13g2_decap_8
XFILLER_9_406 VDD VSS sg13g2_decap_8
XFILLER_22_980 VDD VSS sg13g2_decap_8
XFILLER_43_98 VDD VSS sg13g2_decap_8
XFILLER_40_265 VDD VSS sg13g2_fill_2
XFILLER_40_276 VDD VSS sg13g2_fill_2
XFILLER_21_490 VDD VSS sg13g2_decap_8
XFILLER_5_623 VDD VSS sg13g2_decap_8
XFILLER_111_0 VDD VSS sg13g2_decap_8
XFILLER_4_133 VDD VSS sg13g2_decap_8
XFILLER_107_562 VDD VSS sg13g2_decap_8
XFILLER_49_1042 VDD VSS sg13g2_decap_8
XFILLER_96_906 VDD VSS sg13g2_decap_8
XFILLER_108_91 VDD VSS sg13g2_decap_8
XFILLER_68_608 VDD VSS sg13g2_decap_8
XFILLER_1_840 VDD VSS sg13g2_decap_8
XFILLER_95_427 VDD VSS sg13g2_decap_8
XFILLER_49_811 VDD VSS sg13g2_decap_8
XFILLER_0_350 VDD VSS sg13g2_decap_8
XFILLER_48_343 VDD VSS sg13g2_decap_8
XFILLER_76_685 VDD VSS sg13g2_decap_8
XFILLER_75_140 VDD VSS sg13g2_decap_8
XFILLER_91_644 VDD VSS sg13g2_decap_8
XFILLER_64_858 VDD VSS sg13g2_decap_4
XFILLER_63_324 VDD VSS sg13g2_decap_8
XFILLER_1_1022 VDD VSS sg13g2_decap_8
XFILLER_32_700 VDD VSS sg13g2_decap_8
XFILLER_17_763 VDD VSS sg13g2_decap_8
XFILLER_44_571 VDD VSS sg13g2_decap_8
XFILLER_16_273 VDD VSS sg13g2_decap_8
XFILLER_31_210 VDD VSS sg13g2_decap_8
XFILLER_56_1057 VDD VSS sg13g2_decap_4
XFILLER_17_1008 VDD VSS sg13g2_decap_8
XFILLER_20_917 VDD VSS sg13g2_decap_8
XFILLER_32_777 VDD VSS sg13g2_decap_8
XFILLER_13_980 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_11_clk clkbuf_2_2__f_clk/X clkload8/A VDD VSS sg13g2_buf_8
XFILLER_12_490 VDD VSS sg13g2_decap_8
XFILLER_31_287 VDD VSS sg13g2_decap_8
X_1703_ _1709_/A _1703_/A _1715_/A VDD VSS sg13g2_xnor2_1
XFILLER_9_973 VDD VSS sg13g2_decap_8
XFILLER_8_483 VDD VSS sg13g2_decap_8
XFILLER_99_722 VDD VSS sg13g2_decap_8
X_1634_ _1634_/Y _1634_/A _1634_/B VDD VSS sg13g2_nand2_1
XFILLER_98_232 VDD VSS sg13g2_decap_8
X_2185__170 VDD VSS _2185_/RESET_B sg13g2_tiehi
X_1565_ VSS VDD _1573_/A1 _1210_/Y _1565_/Y _1523_/B sg13g2_a21oi_1
XFILLER_87_917 VDD VSS sg13g2_decap_8
XFILLER_99_766 VDD VSS sg13g2_decap_8
XFILLER_86_405 VDD VSS sg13g2_decap_8
X_1496_ VSS VDD _2266_/Q _1495_/C _1496_/Y _1495_/A sg13g2_a21oi_1
XFILLER_58_107 VDD VSS sg13g2_decap_8
XFILLER_95_994 VDD VSS sg13g2_decap_8
XFILLER_82_611 VDD VSS sg13g2_decap_8
XFILLER_104_49 VDD VSS sg13g2_decap_8
XFILLER_67_663 VDD VSS sg13g2_decap_8
XFILLER_55_825 VDD VSS sg13g2_decap_8
XFILLER_94_482 VDD VSS sg13g2_decap_8
X_2117_ _2117_/Y _2124_/B _2117_/B VDD VSS sg13g2_nand2_1
XFILLER_66_195 VDD VSS sg13g2_decap_8
XFILLER_54_313 VDD VSS sg13g2_decap_8
XFILLER_39_387 VDD VSS sg13g2_decap_8
XFILLER_82_688 VDD VSS sg13g2_decap_8
X_2048_ _2061_/S _2069_/S _2048_/A _2075_/B VDD VSS sg13g2_nand3_1
XFILLER_23_700 VDD VSS sg13g2_decap_8
XFILLER_35_560 VDD VSS sg13g2_decap_8
XFILLER_22_210 VDD VSS sg13g2_decap_8
Xfanout14 _1826_/B _2040_/A VDD VSS sg13g2_buf_1
Xfanout36 fanout40/X _1344_/A2 VDD VSS sg13g2_buf_1
Xfanout47 _2310_/Q _1674_/B VDD VSS sg13g2_buf_1
Xfanout25 _1453_/B _1463_/B VDD VSS sg13g2_buf_1
Xfanout69 _1228_/A _1670_/A VDD VSS sg13g2_buf_1
XFILLER_50_574 VDD VSS sg13g2_decap_8
XFILLER_23_777 VDD VSS sg13g2_decap_8
XFILLER_11_917 VDD VSS sg13g2_decap_8
Xfanout58 _2284_/Q _1634_/A VDD VSS sg13g2_buf_1
XFILLER_109_805 VDD VSS sg13g2_decap_8
XFILLER_10_427 VDD VSS sg13g2_decap_8
XFILLER_13_35 VDD VSS sg13g2_decap_8
XFILLER_22_287 VDD VSS sg13g2_decap_8
XFILLER_108_326 VDD VSS sg13g2_decap_8
XFILLER_89_28 VDD VSS sg13g2_decap_8
Xhold472 _2319_/Q VDD VSS hold472/X sg13g2_dlygate4sd3_1
XFILLER_89_221 VDD VSS sg13g2_decap_4
Xhold450 _2298_/Q VDD VSS _1674_/A sg13g2_dlygate4sd3_1
Xhold461 _2279_/Q VDD VSS hold461/X sg13g2_dlygate4sd3_1
XFILLER_2_637 VDD VSS sg13g2_decap_8
Xhold483 _2222_/Q VDD VSS hold483/X sg13g2_dlygate4sd3_1
XFILLER_89_265 VDD VSS sg13g2_decap_8
Xhold494 _2211_/Q VDD VSS _1368_/A sg13g2_dlygate4sd3_1
XFILLER_77_405 VDD VSS sg13g2_decap_8
XFILLER_1_147 VDD VSS sg13g2_decap_8
XFILLER_104_598 VDD VSS sg13g2_decap_8
XFILLER_38_21 VDD VSS sg13g2_decap_8
XFILLER_58_630 VDD VSS sg13g2_decap_8
XFILLER_86_972 VDD VSS sg13g2_decap_8
XFILLER_73_600 VDD VSS sg13g2_decap_4
XFILLER_46_803 VDD VSS sg13g2_decap_8
XFILLER_79_1024 VDD VSS sg13g2_fill_1
XFILLER_100_793 VDD VSS sg13g2_decap_8
XFILLER_85_482 VDD VSS sg13g2_decap_8
XFILLER_38_98 VDD VSS sg13g2_decap_8
XFILLER_72_154 VDD VSS sg13g2_decap_8
X_2316__246 VDD VSS _2316_/RESET_B sg13g2_tiehi
XFILLER_26_560 VDD VSS sg13g2_decap_8
XFILLER_60_338 VDD VSS sg13g2_decap_8
X_2355__273 VDD VSS _2355_/RESET_B sg13g2_tiehi
XFILLER_14_700 VDD VSS sg13g2_decap_8
XFILLER_54_42 VDD VSS sg13g2_fill_1
XFILLER_54_64 VDD VSS sg13g2_decap_8
XFILLER_13_210 VDD VSS sg13g2_decap_8
XFILLER_110_70 VDD VSS sg13g2_decap_8
XFILLER_9_203 VDD VSS sg13g2_decap_8
XFILLER_14_777 VDD VSS sg13g2_decap_8
XFILLER_13_287 VDD VSS sg13g2_decap_8
XFILLER_103_1022 VDD VSS sg13g2_decap_8
XFILLER_70_63 VDD VSS sg13g2_decap_8
XFILLER_6_910 VDD VSS sg13g2_decap_8
XFILLER_5_420 VDD VSS sg13g2_decap_8
XFILLER_10_994 VDD VSS sg13g2_decap_8
XFILLER_108_871 VDD VSS sg13g2_decap_8
XFILLER_6_987 VDD VSS sg13g2_decap_8
XFILLER_107_370 VDD VSS sg13g2_fill_2
XFILLER_107_381 VDD VSS sg13g2_decap_8
XFILLER_5_497 VDD VSS sg13g2_decap_8
XFILLER_48_7 VDD VSS sg13g2_decap_8
XFILLER_96_714 VDD VSS sg13g2_decap_8
X_1350_ _1351_/A _1347_/Y hold488/X _1347_/B _1370_/A VDD VSS sg13g2_a22oi_1
XFILLER_96_747 VDD VSS sg13g2_decap_8
XFILLER_68_427 VDD VSS sg13g2_decap_8
X_1281_ VDD _2170_/D _1281_/A VSS sg13g2_inv_1
XFILLER_110_557 VDD VSS sg13g2_decap_8
XFILLER_95_257 VDD VSS sg13g2_fill_1
XFILLER_23_1001 VDD VSS sg13g2_decap_8
XFILLER_92_920 VDD VSS sg13g2_fill_2
XFILLER_77_972 VDD VSS sg13g2_decap_8
XFILLER_95_279 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_0_clk clkbuf_leaf_0_clk/A clkload0/A VDD VSS sg13g2_buf_8
XFILLER_110_1026 VDD VSS sg13g2_decap_8
XFILLER_92_953 VDD VSS sg13g2_decap_8
XFILLER_37_847 VDD VSS sg13g2_decap_8
XFILLER_64_655 VDD VSS sg13g2_decap_8
XFILLER_52_817 VDD VSS sg13g2_decap_8
XFILLER_36_357 VDD VSS sg13g2_decap_8
XFILLER_91_496 VDD VSS sg13g2_fill_2
XFILLER_45_891 VDD VSS sg13g2_fill_1
XFILLER_51_305 VDD VSS sg13g2_decap_8
XFILLER_17_560 VDD VSS sg13g2_decap_8
XFILLER_60_872 VDD VSS sg13g2_decap_8
XFILLER_32_574 VDD VSS sg13g2_decap_8
XFILLER_20_714 VDD VSS sg13g2_decap_8
XFILLER_74_0 VDD VSS sg13g2_decap_8
XFILLER_9_770 VDD VSS sg13g2_decap_8
XFILLER_8_280 VDD VSS sg13g2_decap_8
X_1617_ _1623_/A _1617_/A _1629_/A VDD VSS sg13g2_xnor2_1
XFILLER_99_541 VDD VSS sg13g2_decap_8
XFILLER_87_703 VDD VSS sg13g2_decap_8
XFILLER_5_91 VDD VSS sg13g2_decap_8
XFILLER_101_513 VDD VSS sg13g2_decap_8
X_1548_ _1576_/A _1548_/B _2277_/D VDD VSS sg13g2_nor2_1
X_1479_ VSS VDD _1195_/Y _1479_/A2 _2258_/D _1478_/Y sg13g2_a21oi_1
XFILLER_83_920 VDD VSS sg13g2_decap_4
XFILLER_39_140 VDD VSS sg13g2_decap_8
XFILLER_83_953 VDD VSS sg13g2_decap_8
XFILLER_95_780 VDD VSS sg13g2_decap_8
XFILLER_28_847 VDD VSS sg13g2_decap_8
XFILLER_67_471 VDD VSS sg13g2_decap_8
XFILLER_83_986 VDD VSS sg13g2_decap_8
XFILLER_55_655 VDD VSS sg13g2_decap_8
XFILLER_27_357 VDD VSS sg13g2_decap_8
XFILLER_82_485 VDD VSS sg13g2_decap_8
XFILLER_55_699 VDD VSS sg13g2_decap_8
XFILLER_43_828 VDD VSS sg13g2_decap_8
XFILLER_70_647 VDD VSS sg13g2_decap_8
XFILLER_51_883 VDD VSS sg13g2_decap_8
XFILLER_23_574 VDD VSS sg13g2_decap_8
XFILLER_11_714 VDD VSS sg13g2_decap_8
XFILLER_24_56 VDD VSS sg13g2_decap_8
XFILLER_10_224 VDD VSS sg13g2_decap_8
XFILLER_7_707 VDD VSS sg13g2_decap_8
XFILLER_109_602 VDD VSS sg13g2_decap_8
XFILLER_6_217 VDD VSS sg13g2_decap_8
XFILLER_108_112 VDD VSS sg13g2_decap_8
XFILLER_109_679 VDD VSS sg13g2_decap_8
XFILLER_40_77 VDD VSS sg13g2_decap_8
XFILLER_3_924 VDD VSS sg13g2_decap_8
XFILLER_85_1050 VDD VSS sg13g2_decap_8
XFILLER_2_434 VDD VSS sg13g2_decap_8
XFILLER_105_896 VDD VSS sg13g2_decap_8
XFILLER_46_1045 VDD VSS sg13g2_decap_8
XFILLER_49_42 VDD VSS sg13g2_decap_8
XFILLER_104_384 VDD VSS sg13g2_decap_4
XFILLER_77_235 VDD VSS sg13g2_decap_8
XFILLER_59_950 VDD VSS sg13g2_decap_8
XFILLER_93_717 VDD VSS sg13g2_decap_8
XFILLER_92_249 VDD VSS sg13g2_decap_8
XFILLER_105_70 VDD VSS sg13g2_decap_8
XFILLER_1_49 VDD VSS sg13g2_decap_8
XFILLER_19_847 VDD VSS sg13g2_decap_8
XFILLER_73_463 VDD VSS sg13g2_decap_8
XFILLER_18_357 VDD VSS sg13g2_decap_8
XFILLER_45_132 VDD VSS sg13g2_decap_8
XFILLER_65_63 VDD VSS sg13g2_fill_1
XFILLER_61_625 VDD VSS sg13g2_decap_4
XFILLER_60_113 VDD VSS sg13g2_decap_8
XFILLER_42_861 VDD VSS sg13g2_decap_8
XFILLER_60_179 VDD VSS sg13g2_decap_8
XFILLER_14_574 VDD VSS sg13g2_decap_8
XFILLER_81_84 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_10_791 VDD VSS sg13g2_decap_8
XFILLER_6_784 VDD VSS sg13g2_decap_8
X_1402_ VDD _2223_/D _1402_/A VSS sg13g2_inv_1
XFILLER_5_294 VDD VSS sg13g2_decap_8
XFILLER_96_500 VDD VSS sg13g2_decap_8
XFILLER_111_833 VDD VSS sg13g2_decap_8
XFILLER_69_769 VDD VSS sg13g2_decap_8
XFILLER_110_310 VDD VSS sg13g2_fill_1
X_1333_ VDD _2196_/D _1333_/A VSS sg13g2_inv_1
XFILLER_68_246 VDD VSS sg13g2_decap_8
XFILLER_110_354 VDD VSS sg13g2_decap_8
X_1264_ _2359_/Q _2150_/A _1264_/X VDD VSS sg13g2_and2_1
XFILLER_56_419 VDD VSS sg13g2_decap_8
XFILLER_7_1050 VDD VSS sg13g2_decap_8
XFILLER_96_599 VDD VSS sg13g2_decap_8
XFILLER_83_238 VDD VSS sg13g2_decap_4
XFILLER_49_471 VDD VSS sg13g2_decap_8
XFILLER_80_901 VDD VSS sg13g2_decap_8
XFILLER_65_986 VDD VSS sg13g2_decap_8
XFILLER_37_644 VDD VSS sg13g2_decap_8
X_1195_ VDD _1195_/Y _1195_/A VSS sg13g2_inv_1
Xclkbuf_2_1__f_clk clkbuf_leaf_5_clk/A clkbuf_0_clk/X VDD VSS sg13g2_buf_16
XFILLER_52_603 VDD VSS sg13g2_decap_8
XFILLER_36_154 VDD VSS sg13g2_decap_8
XFILLER_101_28 VDD VSS sg13g2_decap_8
XFILLER_40_809 VDD VSS sg13g2_decap_8
XFILLER_33_861 VDD VSS sg13g2_decap_8
XFILLER_51_157 VDD VSS sg13g2_decap_8
XFILLER_20_511 VDD VSS sg13g2_decap_8
XFILLER_32_371 VDD VSS sg13g2_decap_8
XFILLER_20_588 VDD VSS sg13g2_decap_8
XFILLER_105_126 VDD VSS sg13g2_decap_8
XFILLER_10_14 VDD VSS sg13g2_decap_8
XFILLER_102_811 VDD VSS sg13g2_decap_8
XFILLER_99_360 VDD VSS sg13g2_decap_8
XFILLER_87_500 VDD VSS sg13g2_decap_8
XFILLER_0_938 VDD VSS sg13g2_decap_8
XFILLER_87_555 VDD VSS sg13g2_decap_8
XFILLER_102_888 VDD VSS sg13g2_decap_8
XFILLER_75_728 VDD VSS sg13g2_decap_8
XFILLER_101_365 VDD VSS sg13g2_decap_8
XFILLER_19_56 VDD VSS sg13g2_decap_8
XFILLER_47_408 VDD VSS sg13g2_fill_1
XFILLER_74_216 VDD VSS sg13g2_decap_8
XFILLER_28_644 VDD VSS sg13g2_decap_8
XFILLER_55_452 VDD VSS sg13g2_decap_8
XFILLER_83_794 VDD VSS sg13g2_decap_8
XFILLER_82_271 VDD VSS sg13g2_decap_8
XFILLER_70_400 VDD VSS sg13g2_decap_8
XFILLER_43_625 VDD VSS sg13g2_decap_8
XFILLER_27_154 VDD VSS sg13g2_decap_8
XFILLER_71_956 VDD VSS sg13g2_decap_8
XFILLER_70_477 VDD VSS sg13g2_decap_8
XFILLER_24_861 VDD VSS sg13g2_decap_8
XFILLER_35_77 VDD VSS sg13g2_decap_8
XFILLER_30_308 VDD VSS sg13g2_decap_8
XFILLER_11_511 VDD VSS sg13g2_decap_8
XFILLER_51_21 VDD VSS sg13g2_fill_2
XFILLER_23_371 VDD VSS sg13g2_decap_8
XFILLER_7_504 VDD VSS sg13g2_decap_8
XFILLER_11_588 VDD VSS sg13g2_decap_8
XFILLER_13_1022 VDD VSS sg13g2_decap_8
XFILLER_109_476 VDD VSS sg13g2_decap_8
XFILLER_3_721 VDD VSS sg13g2_decap_8
XFILLER_2_231 VDD VSS sg13g2_decap_8
XFILLER_4_0 VDD VSS sg13g2_decap_8
XFILLER_97_308 VDD VSS sg13g2_decap_8
XFILLER_3_798 VDD VSS sg13g2_decap_8
XFILLER_105_693 VDD VSS sg13g2_decap_8
XFILLER_104_181 VDD VSS sg13g2_decap_8
XFILLER_78_522 VDD VSS sg13g2_decap_8
XFILLER_65_205 VDD VSS sg13g2_decap_8
XFILLER_76_84 VDD VSS sg13g2_decap_8
XFILLER_47_931 VDD VSS sg13g2_fill_1
XFILLER_74_750 VDD VSS sg13g2_fill_2
XFILLER_47_964 VDD VSS sg13g2_decap_8
XFILLER_19_644 VDD VSS sg13g2_decap_8
XFILLER_20_1015 VDD VSS sg13g2_decap_8
XFILLER_61_411 VDD VSS sg13g2_decap_8
XFILLER_18_154 VDD VSS sg13g2_decap_8
XFILLER_62_978 VDD VSS sg13g2_fill_1
XFILLER_62_967 VDD VSS sg13g2_decap_8
XFILLER_34_658 VDD VSS sg13g2_decap_8
XFILLER_46_496 VDD VSS sg13g2_decap_8
XFILLER_15_861 VDD VSS sg13g2_decap_8
XFILLER_21_308 VDD VSS sg13g2_decap_8
XFILLER_33_168 VDD VSS sg13g2_decap_8
XFILLER_109_1050 VDD VSS sg13g2_decap_8
X_1951_ _1955_/A _1951_/A _1951_/B VDD VSS sg13g2_xnor2_1
XFILLER_14_371 VDD VSS sg13g2_decap_8
X_1882_ _1887_/A _1887_/B _1882_/Y VDD VSS sg13g2_nor2b_1
XFILLER_30_875 VDD VSS sg13g2_decap_8
XFILLER_6_581 VDD VSS sg13g2_decap_8
XFILLER_111_630 VDD VSS sg13g2_decap_8
XFILLER_97_853 VDD VSS sg13g2_decap_8
XFILLER_69_544 VDD VSS sg13g2_decap_8
X_2365_ _2365_/RESET_B VSS VDD _2365_/D _2365_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_37_0 VDD VSS sg13g2_decap_8
XFILLER_84_503 VDD VSS sg13g2_decap_8
XFILLER_110_140 VDD VSS sg13g2_decap_8
X_1316_ _1316_/Y _1482_/B1 hold389/X _1482_/A2 _2321_/Q VDD VSS sg13g2_a22oi_1
XFILLER_99_1049 VDD VSS sg13g2_decap_8
XFILLER_99_1038 VDD VSS sg13g2_fill_2
XFILLER_96_385 VDD VSS sg13g2_decap_8
XFILLER_2_70 VDD VSS sg13g2_decap_8
X_2296_ _2296_/RESET_B VSS VDD _2296_/D _2296_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_38_975 VDD VSS sg13g2_decap_8
X_2375__232 VDD VSS _2375_/RESET_B sg13g2_tiehi
XFILLER_56_249 VDD VSS sg13g2_decap_8
X_1247_ _1247_/B _1247_/C _1247_/A _1249_/B VDD VSS _1247_/D sg13g2_nand4_1
XFILLER_37_441 VDD VSS sg13g2_decap_8
XFILLER_71_219 VDD VSS sg13g2_decap_8
XFILLER_112_49 VDD VSS sg13g2_decap_8
XFILLER_80_753 VDD VSS sg13g2_decap_8
XFILLER_25_658 VDD VSS sg13g2_decap_8
XFILLER_64_282 VDD VSS sg13g2_decap_8
XFILLER_64_293 VDD VSS sg13g2_decap_8
XFILLER_40_606 VDD VSS sg13g2_decap_8
XFILLER_12_308 VDD VSS sg13g2_decap_8
XFILLER_24_168 VDD VSS sg13g2_decap_8
XFILLER_36_1022 VDD VSS sg13g2_decap_8
XFILLER_52_499 VDD VSS sg13g2_fill_2
XFILLER_52_488 VDD VSS sg13g2_decap_8
XFILLER_21_875 VDD VSS sg13g2_decap_8
X_2312__282 VDD VSS _2312_/RESET_B sg13g2_tiehi
XFILLER_20_385 VDD VSS sg13g2_decap_8
XFILLER_21_35 VDD VSS sg13g2_decap_8
XFILLER_107_947 VDD VSS sg13g2_decap_8
XFILLER_4_518 VDD VSS sg13g2_decap_8
XFILLER_106_435 VDD VSS sg13g2_decap_8
XFILLER_97_28 VDD VSS sg13g2_decap_8
XFILLER_102_630 VDD VSS sg13g2_decap_8
XFILLER_87_330 VDD VSS sg13g2_decap_8
XFILLER_0_735 VDD VSS sg13g2_decap_8
XFILLER_88_886 VDD VSS sg13g2_decap_8
XFILLER_101_140 VDD VSS sg13g2_decap_8
XFILLER_48_717 VDD VSS sg13g2_fill_1
XFILLER_75_514 VDD VSS sg13g2_decap_8
XFILLER_101_151 VDD VSS sg13g2_fill_1
XFILLER_43_1059 VDD VSS sg13g2_fill_2
XFILLER_29_931 VDD VSS sg13g2_decap_8
XFILLER_47_205 VDD VSS sg13g2_decap_8
XFILLER_63_709 VDD VSS sg13g2_decap_8
XFILLER_46_21 VDD VSS sg13g2_decap_8
XFILLER_28_441 VDD VSS sg13g2_decap_8
XFILLER_47_238 VDD VSS sg13g2_decap_8
XFILLER_90_528 VDD VSS sg13g2_decap_8
XFILLER_71_720 VDD VSS sg13g2_decap_8
XFILLER_44_956 VDD VSS sg13g2_decap_8
XFILLER_16_658 VDD VSS sg13g2_decap_8
XFILLER_46_98 VDD VSS sg13g2_decap_4
XFILLER_70_241 VDD VSS sg13g2_decap_8
XFILLER_15_168 VDD VSS sg13g2_decap_8
XFILLER_43_455 VDD VSS sg13g2_decap_8
XFILLER_70_285 VDD VSS sg13g2_decap_8
XFILLER_30_105 VDD VSS sg13g2_decap_8
XFILLER_62_42 VDD VSS sg13g2_decap_8
X_2348__109 VDD VSS _2348_/RESET_B sg13g2_tiehi
XFILLER_7_301 VDD VSS sg13g2_decap_8
XFILLER_12_875 VDD VSS sg13g2_decap_8
XFILLER_109_240 VDD VSS sg13g2_decap_8
XFILLER_11_385 VDD VSS sg13g2_decap_8
XFILLER_8_868 VDD VSS sg13g2_decap_8
XFILLER_7_378 VDD VSS sg13g2_decap_8
XFILLER_98_606 VDD VSS sg13g2_fill_2
XFILLER_97_105 VDD VSS sg13g2_decap_8
XFILLER_79_842 VDD VSS sg13g2_fill_2
XFILLER_112_427 VDD VSS sg13g2_decap_8
XFILLER_105_490 VDD VSS sg13g2_decap_8
XFILLER_3_595 VDD VSS sg13g2_decap_8
XFILLER_30_7 VDD VSS sg13g2_decap_8
XFILLER_39_717 VDD VSS sg13g2_decap_8
XFILLER_78_396 VDD VSS sg13g2_decap_8
X_2150_ _2150_/A _2150_/B _2262_/D VDD VSS sg13g2_and2_1
XFILLER_94_878 VDD VSS sg13g2_decap_8
X_2081_ VSS VDD _2061_/S _2055_/B _2081_/Y _2004_/B sg13g2_a21oi_1
XFILLER_93_355 VDD VSS sg13g2_decap_8
XFILLER_66_547 VDD VSS sg13g2_decap_8
XFILLER_47_750 VDD VSS sg13g2_decap_8
XFILLER_19_441 VDD VSS sg13g2_decap_8
XFILLER_38_238 VDD VSS sg13g2_decap_8
XFILLER_98_1060 VDD VSS sg13g2_fill_1
XFILLER_81_517 VDD VSS sg13g2_decap_8
XFILLER_59_1055 VDD VSS sg13g2_decap_4
XFILLER_35_945 VDD VSS sg13g2_decap_8
XFILLER_62_775 VDD VSS sg13g2_decap_8
XFILLER_50_904 VDD VSS sg13g2_decap_8
XFILLER_61_241 VDD VSS sg13g2_fill_1
X_2290__149 VDD VSS _2290_/RESET_B sg13g2_tiehi
XFILLER_34_455 VDD VSS sg13g2_decap_8
XFILLER_21_105 VDD VSS sg13g2_decap_8
X_1934_ _1935_/A _1934_/A _1934_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_672 VDD VSS sg13g2_decap_8
X_2231__291 VDD VSS _2231_/RESET_B sg13g2_tiehi
X_1865_ _1852_/C _1852_/B _1852_/A _1866_/B VDD VSS sg13g2_a21o_1
X_1796_ _2226_/Q _2218_/Q _1825_/A VDD VSS sg13g2_xor2_1
XFILLER_89_617 VDD VSS sg13g2_decap_8
XFILLER_88_105 VDD VSS sg13g2_decap_8
XFILLER_107_49 VDD VSS sg13g2_decap_8
XFILLER_97_661 VDD VSS sg13g2_decap_8
XFILLER_69_341 VDD VSS sg13g2_decap_8
XFILLER_112_994 VDD VSS sg13g2_decap_8
X_2348_ _2348_/RESET_B VSS VDD _2348_/D _2348_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_57_514 VDD VSS sg13g2_decap_8
XFILLER_96_182 VDD VSS sg13g2_decap_8
XFILLER_84_355 VDD VSS sg13g2_decap_8
X_2279_ _2279_/RESET_B VSS VDD _2279_/D _2279_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_29_238 VDD VSS sg13g2_decap_8
XFILLER_38_772 VDD VSS sg13g2_decap_8
XFILLER_84_399 VDD VSS sg13g2_decap_4
XFILLER_26_945 VDD VSS sg13g2_decap_8
X_2195__150 VDD VSS _2195_/RESET_B sg13g2_tiehi
XFILLER_16_35 VDD VSS sg13g2_decap_8
XFILLER_25_455 VDD VSS sg13g2_decap_8
XFILLER_41_937 VDD VSS sg13g2_decap_8
XFILLER_12_105 VDD VSS sg13g2_decap_8
XFILLER_52_274 VDD VSS sg13g2_decap_8
XFILLER_40_447 VDD VSS sg13g2_decap_8
XFILLER_21_672 VDD VSS sg13g2_decap_8
XFILLER_32_56 VDD VSS sg13g2_decap_8
XFILLER_20_182 VDD VSS sg13g2_decap_8
XFILLER_5_805 VDD VSS sg13g2_decap_8
XFILLER_4_315 VDD VSS sg13g2_decap_8
XFILLER_107_744 VDD VSS sg13g2_decap_8
XFILLER_106_210 VDD VSS sg13g2_decap_8
XFILLER_10_1036 VDD VSS sg13g2_decap_8
XFILLER_79_105 VDD VSS sg13g2_decap_8
XFILLER_106_298 VDD VSS sg13g2_decap_8
XFILLER_88_661 VDD VSS sg13g2_decap_4
XFILLER_0_532 VDD VSS sg13g2_decap_8
XFILLER_103_994 VDD VSS sg13g2_decap_8
XFILLER_88_672 VDD VSS sg13g2_decap_8
XFILLER_76_823 VDD VSS sg13g2_decap_8
XFILLER_94_119 VDD VSS sg13g2_decap_8
XFILLER_48_503 VDD VSS sg13g2_decap_8
XFILLER_75_355 VDD VSS sg13g2_decap_8
XFILLER_91_815 VDD VSS sg13g2_decap_8
XFILLER_91_826 VDD VSS sg13g2_fill_2
XFILLER_63_517 VDD VSS sg13g2_decap_8
XFILLER_90_347 VDD VSS sg13g2_fill_1
XFILLER_17_945 VDD VSS sg13g2_decap_8
XFILLER_71_550 VDD VSS sg13g2_decap_8
XFILLER_73_63 VDD VSS sg13g2_decap_8
XFILLER_44_753 VDD VSS sg13g2_decap_8
XFILLER_16_455 VDD VSS sg13g2_decap_8
XFILLER_32_959 VDD VSS sg13g2_decap_8
XFILLER_19_1050 VDD VSS sg13g2_decap_8
XFILLER_31_469 VDD VSS sg13g2_decap_8
XFILLER_106_1042 VDD VSS sg13g2_decap_8
XFILLER_40_970 VDD VSS sg13g2_decap_8
XFILLER_12_672 VDD VSS sg13g2_decap_8
XFILLER_78_7 VDD VSS sg13g2_decap_8
XFILLER_11_182 VDD VSS sg13g2_decap_8
XFILLER_8_665 VDD VSS sg13g2_decap_8
X_1650_ _1674_/B _2329_/Q _2321_/Q _2344_/Q _2336_/Q _1677_/A _1650_/X VDD VSS sg13g2_mux4_1
XFILLER_7_175 VDD VSS sg13g2_decap_8
X_1581_ _1580_/Y VDD _1581_/Y VSS _2288_/Q _1578_/Y sg13g2_o21ai_1
XFILLER_112_224 VDD VSS sg13g2_decap_8
XFILLER_98_425 VDD VSS sg13g2_decap_8
XFILLER_4_882 VDD VSS sg13g2_decap_8
XFILLER_79_650 VDD VSS sg13g2_decap_8
XFILLER_100_408 VDD VSS sg13g2_decap_4
XFILLER_98_469 VDD VSS sg13g2_decap_8
XFILLER_3_392 VDD VSS sg13g2_decap_8
XFILLER_26_1043 VDD VSS sg13g2_decap_8
XFILLER_67_834 VDD VSS sg13g2_decap_8
X_2202_ _2202_/RESET_B VSS VDD _2202_/D _2202_/Q clkload9/A sg13g2_dfrbpq_1
X_2133_ VDD VSS _2124_/B _2120_/A _2132_/X hold322/X _2135_/A _2124_/Y sg13g2_a221oi_1
XFILLER_66_322 VDD VSS sg13g2_decap_8
XFILLER_39_536 VDD VSS sg13g2_decap_4
XFILLER_96_1019 VDD VSS sg13g2_decap_4
XFILLER_67_889 VDD VSS sg13g2_decap_8
XFILLER_66_355 VDD VSS sg13g2_decap_8
XFILLER_66_366 VDD VSS sg13g2_fill_2
XFILLER_82_848 VDD VSS sg13g2_decap_8
X_2064_ _2050_/X _2063_/X _2079_/S _2065_/C VDD VSS sg13g2_mux2_1
XFILLER_93_185 VDD VSS sg13g2_decap_4
XFILLER_81_347 VDD VSS sg13g2_fill_1
XFILLER_35_742 VDD VSS sg13g2_decap_8
XFILLER_66_399 VDD VSS sg13g2_decap_8
XFILLER_62_561 VDD VSS sg13g2_decap_8
XFILLER_34_252 VDD VSS sg13g2_decap_8
XFILLER_90_881 VDD VSS sg13g2_decap_8
XFILLER_23_959 VDD VSS sg13g2_decap_8
XFILLER_50_756 VDD VSS sg13g2_decap_8
XFILLER_10_609 VDD VSS sg13g2_decap_8
XFILLER_22_469 VDD VSS sg13g2_decap_8
XFILLER_108_508 VDD VSS sg13g2_decap_8
X_1917_ _1919_/B _1917_/A _1917_/B VDD VSS sg13g2_xnor2_1
XFILLER_33_1036 VDD VSS sg13g2_decap_8
X_1848_ VDD _1856_/B _1848_/A VSS sg13g2_inv_1
XFILLER_8_91 VDD VSS sg13g2_decap_8
XFILLER_104_703 VDD VSS sg13g2_decap_8
X_1779_ _2213_/Q _2221_/Q _1779_/Y VDD VSS sg13g2_nor2b_1
XFILLER_2_819 VDD VSS sg13g2_decap_8
XFILLER_104_736 VDD VSS sg13g2_decap_8
XFILLER_1_329 VDD VSS sg13g2_decap_8
XFILLER_103_235 VDD VSS sg13g2_decap_8
XFILLER_76_119 VDD VSS sg13g2_decap_8
XFILLER_112_791 VDD VSS sg13g2_decap_8
XFILLER_85_631 VDD VSS sg13g2_fill_2
XFILLER_85_642 VDD VSS sg13g2_fill_2
XFILLER_85_675 VDD VSS sg13g2_decap_8
XFILLER_84_163 VDD VSS sg13g2_decap_8
XFILLER_27_56 VDD VSS sg13g2_decap_8
XFILLER_45_539 VDD VSS sg13g2_decap_8
XFILLER_26_742 VDD VSS sg13g2_decap_8
XFILLER_41_734 VDD VSS sg13g2_decap_8
XFILLER_25_252 VDD VSS sg13g2_decap_8
XFILLER_14_959 VDD VSS sg13g2_decap_8
XFILLER_13_469 VDD VSS sg13g2_decap_8
XFILLER_43_77 VDD VSS sg13g2_decap_8
XFILLER_5_602 VDD VSS sg13g2_decap_8
XFILLER_4_112 VDD VSS sg13g2_decap_8
XFILLER_107_541 VDD VSS sg13g2_decap_8
XFILLER_104_0 VDD VSS sg13g2_decap_8
XFILLER_5_679 VDD VSS sg13g2_decap_8
XFILLER_108_70 VDD VSS sg13g2_decap_8
XFILLER_4_189 VDD VSS sg13g2_decap_8
XFILLER_4_49 VDD VSS sg13g2_decap_8
XFILLER_95_406 VDD VSS sg13g2_decap_8
XFILLER_110_739 VDD VSS sg13g2_decap_8
XFILLER_1_896 VDD VSS sg13g2_decap_8
XFILLER_67_119 VDD VSS sg13g2_decap_8
XFILLER_68_96 VDD VSS sg13g2_decap_8
XFILLER_103_791 VDD VSS sg13g2_decap_8
XFILLER_49_867 VDD VSS sg13g2_fill_1
XFILLER_49_856 VDD VSS sg13g2_decap_8
XFILLER_48_322 VDD VSS sg13g2_decap_8
XFILLER_76_664 VDD VSS sg13g2_decap_8
XFILLER_91_623 VDD VSS sg13g2_decap_8
XFILLER_75_185 VDD VSS sg13g2_decap_8
XFILLER_90_122 VDD VSS sg13g2_decap_8
XFILLER_64_837 VDD VSS sg13g2_decap_8
XFILLER_1_1001 VDD VSS sg13g2_decap_8
XFILLER_36_539 VDD VSS sg13g2_decap_8
XFILLER_48_388 VDD VSS sg13g2_decap_8
XFILLER_84_84 VDD VSS sg13g2_decap_8
XFILLER_44_550 VDD VSS sg13g2_decap_8
XFILLER_17_742 VDD VSS sg13g2_decap_8
XFILLER_90_188 VDD VSS sg13g2_decap_8
XFILLER_56_1036 VDD VSS sg13g2_decap_8
XFILLER_16_252 VDD VSS sg13g2_decap_8
XFILLER_32_756 VDD VSS sg13g2_decap_8
XFILLER_31_266 VDD VSS sg13g2_decap_8
XFILLER_9_952 VDD VSS sg13g2_decap_8
X_1702_ _1715_/A _2316_/Q _2302_/Q VDD VSS sg13g2_xnor2_1
X_2225__90 VDD VSS _2225__90/L_HI sg13g2_tiehi
XFILLER_8_462 VDD VSS sg13g2_decap_8
X_1633_ _1634_/B _1633_/A _1633_/B VDD VSS sg13g2_xnor2_1
XFILLER_99_701 VDD VSS sg13g2_decap_8
XFILLER_98_211 VDD VSS sg13g2_decap_8
X_1564_ VDD _1564_/Y _1564_/A VSS sg13g2_inv_1
XFILLER_101_706 VDD VSS sg13g2_decap_8
XFILLER_63_1029 VDD VSS sg13g2_fill_1
XIO_FILL_IO_EAST_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_59_609 VDD VSS sg13g2_decap_8
X_1495_ _1497_/B _1495_/A _2266_/Q _1495_/C VDD VSS sg13g2_and3_1
XFILLER_67_642 VDD VSS sg13g2_decap_8
XFILLER_95_973 VDD VSS sg13g2_decap_8
XFILLER_94_461 VDD VSS sg13g2_decap_8
XFILLER_104_28 VDD VSS sg13g2_decap_8
XFILLER_55_804 VDD VSS sg13g2_decap_8
XFILLER_39_366 VDD VSS sg13g2_decap_8
X_2116_ _2144_/S0 hold314/X hold389/X hold308/X hold336/X _1510_/B _2117_/B VDD VSS
+ sg13g2_mux4_1
XFILLER_66_174 VDD VSS sg13g2_decap_8
XFILLER_27_539 VDD VSS sg13g2_decap_8
XFILLER_82_667 VDD VSS sg13g2_decap_8
X_2047_ _2048_/A _2069_/S _2047_/X VDD VSS sg13g2_and2_1
XFILLER_70_829 VDD VSS sg13g2_decap_8
XFILLER_63_881 VDD VSS sg13g2_decap_8
Xfanout15 _1825_/Y _1826_/B VDD VSS sg13g2_buf_1
Xfanout26 _1453_/B _1455_/B VDD VSS sg13g2_buf_1
Xfanout37 fanout40/X _1280_/A2 VDD VSS sg13g2_buf_1
XFILLER_23_756 VDD VSS sg13g2_decap_8
Xfanout48 _1724_/S _1720_/A VDD VSS sg13g2_buf_1
Xfanout59 _2144_/S1 _1510_/B VDD VSS sg13g2_buf_1
XFILLER_50_553 VDD VSS sg13g2_decap_8
XFILLER_10_406 VDD VSS sg13g2_decap_8
XFILLER_13_14 VDD VSS sg13g2_decap_8
XFILLER_22_266 VDD VSS sg13g2_decap_8
XFILLER_50_597 VDD VSS sg13g2_decap_8
XFILLER_108_305 VDD VSS sg13g2_decap_8
XFILLER_89_200 VDD VSS sg13g2_decap_8
Xhold451 _1675_/Y VDD VSS _2310_/D sg13g2_dlygate4sd3_1
XFILLER_8_7 VDD VSS sg13g2_decap_8
XFILLER_2_616 VDD VSS sg13g2_decap_8
Xhold440 _1595_/Y VDD VSS _2289_/D sg13g2_dlygate4sd3_1
Xhold462 _1561_/Y VDD VSS _1562_/B sg13g2_dlygate4sd3_1
Xhold473 _1721_/Y VDD VSS _1722_/B sg13g2_dlygate4sd3_1
Xhold495 _2225_/Q VDD VSS hold495/X sg13g2_dlygate4sd3_1
XFILLER_89_244 VDD VSS sg13g2_decap_8
XFILLER_1_126 VDD VSS sg13g2_decap_8
Xhold484 _2281_/Q VDD VSS hold484/X sg13g2_dlygate4sd3_1
XFILLER_104_577 VDD VSS sg13g2_decap_8
XFILLER_86_951 VDD VSS sg13g2_decap_8
XFILLER_100_772 VDD VSS sg13g2_decap_8
XFILLER_100_750 VDD VSS sg13g2_decap_4
X_2201__138 VDD VSS _2201_/RESET_B sg13g2_tiehi
XFILLER_85_461 VDD VSS sg13g2_decap_4
XFILLER_58_686 VDD VSS sg13g2_decap_8
XFILLER_38_77 VDD VSS sg13g2_decap_8
XFILLER_73_623 VDD VSS sg13g2_decap_8
XFILLER_18_539 VDD VSS sg13g2_decap_8
XFILLER_45_336 VDD VSS sg13g2_decap_8
XFILLER_61_818 VDD VSS sg13g2_decap_4
XFILLER_54_21 VDD VSS sg13g2_fill_2
XFILLER_54_892 VDD VSS sg13g2_decap_8
XFILLER_14_756 VDD VSS sg13g2_decap_8
XFILLER_13_266 VDD VSS sg13g2_decap_8
XFILLER_103_1001 VDD VSS sg13g2_decap_8
XFILLER_70_42 VDD VSS sg13g2_decap_8
XFILLER_9_259 VDD VSS sg13g2_decap_8
XFILLER_10_973 VDD VSS sg13g2_decap_8
XFILLER_108_850 VDD VSS sg13g2_decap_8
XFILLER_6_966 VDD VSS sg13g2_decap_8
XFILLER_107_360 VDD VSS sg13g2_decap_8
XFILLER_5_476 VDD VSS sg13g2_decap_8
XFILLER_79_84 VDD VSS sg13g2_decap_8
XFILLER_69_929 VDD VSS sg13g2_decap_8
XFILLER_95_203 VDD VSS sg13g2_decap_4
XFILLER_68_406 VDD VSS sg13g2_decap_8
XFILLER_77_951 VDD VSS sg13g2_decap_8
X_1280_ _1280_/Y _1280_/B1 hold312/X _1280_/A2 _2320_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_536 VDD VSS sg13g2_decap_8
XFILLER_1_693 VDD VSS sg13g2_decap_8
XFILLER_37_826 VDD VSS sg13g2_decap_8
XFILLER_110_1005 VDD VSS sg13g2_decap_8
XFILLER_92_932 VDD VSS sg13g2_decap_8
XFILLER_76_483 VDD VSS sg13g2_decap_8
XFILLER_23_1057 VDD VSS sg13g2_decap_4
XFILLER_64_634 VDD VSS sg13g2_decap_8
XFILLER_49_697 VDD VSS sg13g2_decap_8
XFILLER_63_111 VDD VSS sg13g2_decap_8
XFILLER_36_336 VDD VSS sg13g2_decap_8
XFILLER_48_196 VDD VSS sg13g2_decap_8
XFILLER_91_475 VDD VSS sg13g2_decap_8
XFILLER_63_166 VDD VSS sg13g2_decap_8
XFILLER_60_851 VDD VSS sg13g2_decap_8
XFILLER_63_199 VDD VSS sg13g2_decap_4
XFILLER_32_553 VDD VSS sg13g2_decap_8
XFILLER_67_0 VDD VSS sg13g2_decap_8
XFILLER_99_520 VDD VSS sg13g2_decap_8
X_1616_ _1629_/A _2293_/Q _2278_/Q VDD VSS sg13g2_xnor2_1
XFILLER_5_70 VDD VSS sg13g2_decap_8
XFILLER_99_597 VDD VSS sg13g2_decap_8
XFILLER_86_203 VDD VSS sg13g2_fill_2
X_1547_ _1547_/Y _1527_/Y _1546_/Y hold457/X _1527_/B VDD VSS sg13g2_a22oi_1
XFILLER_8_1029 VDD VSS sg13g2_decap_8
XFILLER_87_759 VDD VSS sg13g2_decap_8
X_1478_ _1602_/B VDD _1478_/Y VSS _1385_/A _1481_/A2 sg13g2_o21ai_1
XFILLER_86_258 VDD VSS sg13g2_decap_8
XFILLER_68_984 VDD VSS sg13g2_decap_4
XFILLER_68_962 VDD VSS sg13g2_decap_4
XFILLER_67_450 VDD VSS sg13g2_decap_8
XFILLER_55_634 VDD VSS sg13g2_decap_8
XFILLER_28_826 VDD VSS sg13g2_decap_8
XFILLER_43_807 VDD VSS sg13g2_decap_8
XFILLER_27_336 VDD VSS sg13g2_decap_8
XFILLER_39_196 VDD VSS sg13g2_decap_8
XFILLER_70_626 VDD VSS sg13g2_decap_8
XFILLER_82_464 VDD VSS sg13g2_decap_8
XFILLER_39_1053 VDD VSS sg13g2_decap_8
XFILLER_23_553 VDD VSS sg13g2_decap_8
XFILLER_24_35 VDD VSS sg13g2_decap_8
XFILLER_10_203 VDD VSS sg13g2_decap_8
XFILLER_109_658 VDD VSS sg13g2_decap_8
XFILLER_108_168 VDD VSS sg13g2_decap_8
XFILLER_3_903 VDD VSS sg13g2_decap_8
XFILLER_40_56 VDD VSS sg13g2_decap_8
XFILLER_108_179 VDD VSS sg13g2_fill_1
XFILLER_2_413 VDD VSS sg13g2_decap_8
XFILLER_78_704 VDD VSS sg13g2_decap_8
XFILLER_46_1024 VDD VSS sg13g2_decap_8
XFILLER_49_21 VDD VSS sg13g2_decap_8
XFILLER_105_875 VDD VSS sg13g2_decap_8
XFILLER_104_363 VDD VSS sg13g2_decap_8
XFILLER_77_203 VDD VSS sg13g2_decap_8
Xhold292 _2363_/Q VDD VSS _1502_/D sg13g2_dlygate4sd3_1
XFILLER_58_450 VDD VSS sg13g2_fill_2
XFILLER_1_28 VDD VSS sg13g2_decap_8
XFILLER_86_781 VDD VSS sg13g2_decap_8
XFILLER_92_228 VDD VSS sg13g2_decap_8
XFILLER_85_280 VDD VSS sg13g2_decap_4
XFILLER_58_483 VDD VSS sg13g2_decap_8
XFILLER_19_826 VDD VSS sg13g2_decap_8
XFILLER_65_42 VDD VSS sg13g2_decap_8
XFILLER_74_954 VDD VSS sg13g2_decap_8
XFILLER_46_645 VDD VSS sg13g2_decap_8
XFILLER_18_336 VDD VSS sg13g2_decap_8
XFILLER_61_637 VDD VSS sg13g2_fill_2
XFILLER_61_604 VDD VSS sg13g2_decap_8
XFILLER_46_689 VDD VSS sg13g2_decap_8
XFILLER_42_840 VDD VSS sg13g2_decap_8
XFILLER_81_63 VDD VSS sg13g2_decap_8
XFILLER_14_553 VDD VSS sg13g2_decap_8
XFILLER_60_147 VDD VSS sg13g2_decap_8
XFILLER_41_350 VDD VSS sg13g2_decap_4
XFILLER_10_770 VDD VSS sg13g2_decap_8
XFILLER_6_763 VDD VSS sg13g2_decap_8
XFILLER_60_7 VDD VSS sg13g2_decap_8
X_2286__165 VDD VSS _2286_/RESET_B sg13g2_tiehi
XFILLER_5_273 VDD VSS sg13g2_decap_8
X_1401_ _1402_/A _1392_/Y hold456/X _1392_/B _1379_/A VDD VSS sg13g2_a22oi_1
XFILLER_111_812 VDD VSS sg13g2_decap_8
XFILLER_69_748 VDD VSS sg13g2_decap_8
XFILLER_110_333 VDD VSS sg13g2_decap_8
X_1332_ _1332_/Y _1344_/B1 hold314/X _1344_/A2 _2329_/Q VDD VSS sg13g2_a22oi_1
XFILLER_68_225 VDD VSS sg13g2_decap_8
XFILLER_2_980 VDD VSS sg13g2_decap_8
XFILLER_111_889 VDD VSS sg13g2_decap_8
XFILLER_96_578 VDD VSS sg13g2_decap_8
XFILLER_83_206 VDD VSS sg13g2_decap_4
X_1263_ _1262_/X hold569/X _1261_/Y _2355_/D VDD VSS sg13g2_a21o_1
XFILLER_1_490 VDD VSS sg13g2_decap_8
XFILLER_77_781 VDD VSS sg13g2_decap_8
XFILLER_37_623 VDD VSS sg13g2_decap_8
XFILLER_49_461 VDD VSS sg13g2_decap_8
XFILLER_65_965 VDD VSS sg13g2_decap_8
XFILLER_36_133 VDD VSS sg13g2_decap_8
X_1194_ VDD _1194_/Y _1194_/A VSS sg13g2_inv_1
XFILLER_92_784 VDD VSS sg13g2_decap_8
XFILLER_64_486 VDD VSS sg13g2_decap_8
XFILLER_33_840 VDD VSS sg13g2_decap_8
XFILLER_32_350 VDD VSS sg13g2_decap_8
XFILLER_20_567 VDD VSS sg13g2_decap_8
XFILLER_69_1024 VDD VSS sg13g2_fill_1
XFILLER_69_1013 VDD VSS sg13g2_fill_1
XFILLER_105_105 VDD VSS sg13g2_decap_8
XFILLER_0_917 VDD VSS sg13g2_decap_8
XFILLER_99_394 VDD VSS sg13g2_fill_2
XFILLER_59_236 VDD VSS sg13g2_decap_8
XFILLER_102_867 VDD VSS sg13g2_decap_8
XFILLER_75_707 VDD VSS sg13g2_decap_8
X_2241__260 VDD VSS _2241_/RESET_B sg13g2_tiehi
XFILLER_101_344 VDD VSS sg13g2_decap_8
XFILLER_19_35 VDD VSS sg13g2_decap_8
XFILLER_28_623 VDD VSS sg13g2_decap_8
XFILLER_83_740 VDD VSS sg13g2_decap_8
XFILLER_67_280 VDD VSS sg13g2_decap_8
XFILLER_55_431 VDD VSS sg13g2_decap_8
XFILLER_27_133 VDD VSS sg13g2_decap_8
XFILLER_76_1028 VDD VSS sg13g2_fill_2
XFILLER_71_935 VDD VSS sg13g2_decap_8
XFILLER_83_773 VDD VSS sg13g2_decap_8
XFILLER_82_250 VDD VSS sg13g2_decap_8
XFILLER_43_604 VDD VSS sg13g2_decap_8
XFILLER_24_840 VDD VSS sg13g2_decap_8
XFILLER_35_56 VDD VSS sg13g2_decap_8
XFILLER_70_456 VDD VSS sg13g2_decap_8
XFILLER_42_147 VDD VSS sg13g2_decap_4
XFILLER_23_350 VDD VSS sg13g2_decap_8
XFILLER_11_567 VDD VSS sg13g2_decap_8
XFILLER_13_1001 VDD VSS sg13g2_decap_8
XFILLER_51_88 VDD VSS sg13g2_decap_8
XFILLER_100_1004 VDD VSS sg13g2_decap_8
XFILLER_109_455 VDD VSS sg13g2_decap_8
XFILLER_100_1059 VDD VSS sg13g2_fill_2
XFILLER_3_700 VDD VSS sg13g2_decap_8
XFILLER_2_210 VDD VSS sg13g2_decap_8
XFILLER_112_609 VDD VSS sg13g2_decap_8
XFILLER_105_672 VDD VSS sg13g2_decap_8
XFILLER_3_777 VDD VSS sg13g2_decap_8
XFILLER_111_119 VDD VSS sg13g2_decap_8
XFILLER_2_287 VDD VSS sg13g2_decap_8
XFILLER_78_578 VDD VSS sg13g2_decap_8
XFILLER_66_707 VDD VSS sg13g2_decap_8
XFILLER_66_729 VDD VSS sg13g2_fill_1
XFILLER_93_526 VDD VSS sg13g2_decap_4
XFILLER_76_63 VDD VSS sg13g2_decap_8
XFILLER_59_770 VDD VSS sg13g2_fill_2
XFILLER_19_623 VDD VSS sg13g2_decap_8
XFILLER_93_548 VDD VSS sg13g2_fill_2
XFILLER_74_740 VDD VSS sg13g2_fill_1
XFILLER_47_943 VDD VSS sg13g2_decap_8
XFILLER_18_133 VDD VSS sg13g2_decap_8
XFILLER_73_250 VDD VSS sg13g2_decap_8
XFILLER_46_453 VDD VSS sg13g2_decap_8
XFILLER_46_475 VDD VSS sg13g2_decap_8
XFILLER_62_946 VDD VSS sg13g2_decap_8
XFILLER_34_637 VDD VSS sg13g2_decap_8
XFILLER_15_840 VDD VSS sg13g2_decap_8
XFILLER_92_84 VDD VSS sg13g2_decap_8
XFILLER_61_467 VDD VSS sg13g2_decap_8
XFILLER_14_350 VDD VSS sg13g2_decap_8
XFILLER_33_147 VDD VSS sg13g2_decap_8
XFILLER_70_990 VDD VSS sg13g2_decap_8
X_1950_ _1950_/Y _1951_/A _1951_/B VDD VSS sg13g2_nand2_1
X_1881_ _1880_/B _1880_/Y _1954_/S _1887_/B VDD VSS sg13g2_mux2_1
XFILLER_30_854 VDD VSS sg13g2_decap_8
XFILLER_6_560 VDD VSS sg13g2_decap_8
XFILLER_103_609 VDD VSS sg13g2_decap_8
XFILLER_69_501 VDD VSS sg13g2_decap_8
XFILLER_97_832 VDD VSS sg13g2_decap_8
XFILLER_102_119 VDD VSS sg13g2_decap_8
X_2364_ _2364_/RESET_B VSS VDD _2364_/D _2364_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_96_364 VDD VSS sg13g2_decap_8
X_1315_ VDD _2187_/D _1315_/A VSS sg13g2_inv_1
XFILLER_111_686 VDD VSS sg13g2_decap_8
XFILLER_84_537 VDD VSS sg13g2_decap_8
X_2295_ _2295_/RESET_B VSS VDD _2295_/D _2295_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_110_196 VDD VSS sg13g2_decap_8
XFILLER_38_954 VDD VSS sg13g2_decap_8
X_1246_ _1248_/C _2292_/Q _2254_/Q VDD VSS sg13g2_xnor2_1
XFILLER_37_420 VDD VSS sg13g2_decap_8
XFILLER_112_28 VDD VSS sg13g2_decap_8
XFILLER_65_773 VDD VSS sg13g2_decap_8
XFILLER_64_261 VDD VSS sg13g2_decap_8
XFILLER_80_732 VDD VSS sg13g2_decap_8
XFILLER_25_637 VDD VSS sg13g2_decap_8
XFILLER_37_497 VDD VSS sg13g2_decap_8
XFILLER_36_1001 VDD VSS sg13g2_decap_8
XFILLER_52_445 VDD VSS sg13g2_decap_8
XFILLER_24_147 VDD VSS sg13g2_decap_8
XFILLER_21_854 VDD VSS sg13g2_decap_8
XFILLER_20_364 VDD VSS sg13g2_decap_8
XFILLER_21_14 VDD VSS sg13g2_decap_8
XFILLER_107_926 VDD VSS sg13g2_decap_8
XFILLER_106_414 VDD VSS sg13g2_decap_8
XFILLER_108_7 VDD VSS sg13g2_decap_8
XFILLER_0_714 VDD VSS sg13g2_decap_8
XFILLER_82_1054 VDD VSS sg13g2_decap_8
XFILLER_88_865 VDD VSS sg13g2_decap_8
XFILLER_99_191 VDD VSS sg13g2_decap_8
XFILLER_43_1038 VDD VSS sg13g2_decap_8
XFILLER_29_910 VDD VSS sg13g2_decap_8
XFILLER_47_217 VDD VSS sg13g2_decap_8
XFILLER_28_420 VDD VSS sg13g2_decap_8
XFILLER_90_518 VDD VSS sg13g2_decap_4
XFILLER_29_987 VDD VSS sg13g2_decap_8
XFILLER_56_784 VDD VSS sg13g2_decap_8
XFILLER_46_77 VDD VSS sg13g2_decap_8
XFILLER_83_592 VDD VSS sg13g2_decap_4
XFILLER_44_935 VDD VSS sg13g2_decap_8
XFILLER_55_294 VDD VSS sg13g2_decap_8
XFILLER_16_637 VDD VSS sg13g2_decap_8
XFILLER_28_497 VDD VSS sg13g2_decap_8
XFILLER_43_434 VDD VSS sg13g2_decap_8
XFILLER_15_147 VDD VSS sg13g2_decap_8
XFILLER_62_21 VDD VSS sg13g2_decap_8
XFILLER_71_798 VDD VSS sg13g2_decap_8
XFILLER_52_990 VDD VSS sg13g2_decap_8
XFILLER_12_854 VDD VSS sg13g2_decap_8
XFILLER_62_98 VDD VSS sg13g2_decap_8
XFILLER_11_364 VDD VSS sg13g2_decap_8
XFILLER_8_847 VDD VSS sg13g2_decap_8
XFILLER_7_357 VDD VSS sg13g2_decap_8
XFILLER_7_49 VDD VSS sg13g2_decap_8
XFILLER_109_263 VDD VSS sg13g2_fill_1
XFILLER_112_406 VDD VSS sg13g2_decap_8
XFILLER_11_91 VDD VSS sg13g2_decap_8
XFILLER_79_821 VDD VSS sg13g2_decap_8
XFILLER_3_574 VDD VSS sg13g2_decap_8
XFILLER_78_342 VDD VSS sg13g2_decap_8
XFILLER_78_353 VDD VSS sg13g2_fill_2
XFILLER_87_84 VDD VSS sg13g2_decap_8
XFILLER_23_7 VDD VSS sg13g2_decap_8
XFILLER_78_375 VDD VSS sg13g2_decap_8
XFILLER_66_526 VDD VSS sg13g2_decap_8
XFILLER_38_217 VDD VSS sg13g2_decap_8
X_2080_ _2080_/Y _2149_/A _2080_/B VDD VSS sg13g2_nand2_1
XFILLER_19_420 VDD VSS sg13g2_decap_8
XFILLER_4_1043 VDD VSS sg13g2_decap_8
XFILLER_35_924 VDD VSS sg13g2_decap_8
XFILLER_74_581 VDD VSS sg13g2_decap_8
XFILLER_59_1034 VDD VSS sg13g2_decap_8
XFILLER_61_220 VDD VSS sg13g2_decap_8
XFILLER_19_497 VDD VSS sg13g2_decap_8
XFILLER_34_434 VDD VSS sg13g2_decap_8
XFILLER_62_754 VDD VSS sg13g2_decap_8
X_1933_ _1938_/A _1933_/A _1933_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_651 VDD VSS sg13g2_decap_8
X_1864_ _1892_/A _1892_/B _1880_/A VDD VSS sg13g2_nor2_1
XIO_FILL_IO_SOUTH_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_1795_ _1795_/A _1801_/B _1811_/A VDD VSS sg13g2_and2_1
XFILLER_104_929 VDD VSS sg13g2_decap_8
XFILLER_107_28 VDD VSS sg13g2_decap_8
XFILLER_66_1049 VDD VSS sg13g2_decap_8
XFILLER_97_640 VDD VSS sg13g2_decap_8
XFILLER_112_973 VDD VSS sg13g2_decap_8
X_2347_ _2347_/RESET_B VSS VDD _2347_/D _2347_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_85_824 VDD VSS sg13g2_decap_8
XFILLER_69_386 VDD VSS sg13g2_decap_8
XFILLER_96_161 VDD VSS sg13g2_decap_8
XFILLER_29_217 VDD VSS sg13g2_decap_8
XFILLER_111_483 VDD VSS sg13g2_decap_8
XFILLER_84_334 VDD VSS sg13g2_decap_8
XFILLER_57_537 VDD VSS sg13g2_fill_1
X_2278_ _2278_/RESET_B VSS VDD _2278_/D _2278_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_72_529 VDD VSS sg13g2_decap_8
XFILLER_26_924 VDD VSS sg13g2_decap_8
XFILLER_38_751 VDD VSS sg13g2_decap_8
X_1229_ _1492_/A _2265_/Q _1465_/B VDD VSS sg13g2_nor2_1
XFILLER_16_14 VDD VSS sg13g2_decap_8
XFILLER_25_434 VDD VSS sg13g2_decap_8
XFILLER_37_294 VDD VSS sg13g2_decap_8
XFILLER_73_1009 VDD VSS sg13g2_decap_8
XFILLER_80_551 VDD VSS sg13g2_decap_8
XFILLER_41_916 VDD VSS sg13g2_decap_8
XFILLER_53_754 VDD VSS sg13g2_decap_8
XFILLER_80_584 VDD VSS sg13g2_decap_8
XFILLER_40_426 VDD VSS sg13g2_decap_8
XFILLER_21_651 VDD VSS sg13g2_decap_8
XFILLER_32_35 VDD VSS sg13g2_decap_8
XFILLER_20_161 VDD VSS sg13g2_decap_8
XFILLER_107_723 VDD VSS sg13g2_decap_8
XFILLER_10_1015 VDD VSS sg13g2_decap_8
XFILLER_106_266 VDD VSS sg13g2_decap_8
XFILLER_0_511 VDD VSS sg13g2_decap_8
XFILLER_88_651 VDD VSS sg13g2_fill_1
XFILLER_103_973 VDD VSS sg13g2_decap_8
XFILLER_87_172 VDD VSS sg13g2_decap_8
XFILLER_0_588 VDD VSS sg13g2_decap_8
XFILLER_57_21 VDD VSS sg13g2_decap_8
XFILLER_57_43 VDD VSS sg13g2_fill_2
XFILLER_87_183 VDD VSS sg13g2_fill_2
XFILLER_75_334 VDD VSS sg13g2_decap_8
XFILLER_48_548 VDD VSS sg13g2_decap_4
XFILLER_76_879 VDD VSS sg13g2_decap_8
X_2319__234 VDD VSS _2319_/RESET_B sg13g2_tiehi
XFILLER_90_326 VDD VSS sg13g2_decap_8
XFILLER_56_581 VDD VSS sg13g2_decap_8
XFILLER_44_732 VDD VSS sg13g2_decap_8
XFILLER_29_784 VDD VSS sg13g2_decap_8
XFILLER_17_924 VDD VSS sg13g2_decap_8
XFILLER_73_42 VDD VSS sg13g2_decap_8
XFILLER_16_434 VDD VSS sg13g2_decap_8
XFILLER_28_294 VDD VSS sg13g2_decap_8
XFILLER_71_573 VDD VSS sg13g2_fill_1
XFILLER_71_584 VDD VSS sg13g2_decap_8
XFILLER_32_938 VDD VSS sg13g2_decap_8
XFILLER_31_448 VDD VSS sg13g2_decap_8
XFILLER_106_1021 VDD VSS sg13g2_decap_8
X_2211__118 VDD VSS _2211_/RESET_B sg13g2_tiehi
XFILLER_12_651 VDD VSS sg13g2_decap_8
XFILLER_11_161 VDD VSS sg13g2_decap_8
XFILLER_8_644 VDD VSS sg13g2_decap_8
XFILLER_7_154 VDD VSS sg13g2_decap_8
X_1580_ _1579_/Y VDD _1580_/Y VSS _1580_/A1 hold449/X sg13g2_o21ai_1
XFILLER_99_938 VDD VSS sg13g2_decap_8
XFILLER_99_927 VDD VSS sg13g2_fill_2
XFILLER_98_404 VDD VSS sg13g2_decap_8
XFILLER_4_861 VDD VSS sg13g2_decap_8
XFILLER_112_203 VDD VSS sg13g2_decap_8
XFILLER_98_448 VDD VSS sg13g2_fill_1
XFILLER_3_371 VDD VSS sg13g2_decap_8
XFILLER_26_1022 VDD VSS sg13g2_decap_8
X_2201_ _2201_/RESET_B VSS VDD _2201_/D _2201_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_66_301 VDD VSS sg13g2_decap_8
X_2132_ _2124_/A _2199_/Q _2191_/Q _2183_/Q _2175_/Q _2144_/S1 _2132_/X VDD VSS sg13g2_mux4_1
XFILLER_94_676 VDD VSS sg13g2_decap_8
XFILLER_94_687 VDD VSS sg13g2_fill_1
XFILLER_82_827 VDD VSS sg13g2_decap_8
XFILLER_67_879 VDD VSS sg13g2_fill_1
XFILLER_66_378 VDD VSS sg13g2_decap_8
XFILLER_75_890 VDD VSS sg13g2_decap_8
X_2063_ _1892_/X _1880_/Y _2069_/S _2063_/X VDD VSS sg13g2_mux2_1
XFILLER_81_326 VDD VSS sg13g2_decap_8
XFILLER_35_721 VDD VSS sg13g2_decap_8
XFILLER_62_540 VDD VSS sg13g2_decap_8
XFILLER_19_294 VDD VSS sg13g2_decap_8
XFILLER_34_231 VDD VSS sg13g2_decap_8
XFILLER_23_938 VDD VSS sg13g2_decap_8
XFILLER_35_798 VDD VSS sg13g2_decap_8
XFILLER_97_0 VDD VSS sg13g2_decap_8
XFILLER_22_448 VDD VSS sg13g2_decap_8
XFILLER_72_1053 VDD VSS sg13g2_decap_8
XFILLER_33_1015 VDD VSS sg13g2_decap_8
X_1916_ _1770_/A VDD _1917_/B VSS _1766_/B _1899_/B sg13g2_o21ai_1
X_1847_ _1848_/A _2248_/Q _2207_/Q VDD VSS sg13g2_xnor2_1
XFILLER_8_70 VDD VSS sg13g2_decap_8
X_1778_ _2214_/Q _2222_/Q _1778_/Y VDD VSS sg13g2_nor2b_1
XFILLER_103_203 VDD VSS sg13g2_decap_4
XFILLER_89_426 VDD VSS sg13g2_decap_8
XFILLER_1_308 VDD VSS sg13g2_decap_8
XFILLER_112_770 VDD VSS sg13g2_decap_8
XFILLER_85_610 VDD VSS sg13g2_decap_8
XFILLER_69_150 VDD VSS sg13g2_fill_1
XFILLER_58_802 VDD VSS sg13g2_decap_8
XFILLER_85_654 VDD VSS sg13g2_decap_8
XFILLER_111_280 VDD VSS sg13g2_decap_8
XFILLER_97_492 VDD VSS sg13g2_fill_2
XFILLER_97_481 VDD VSS sg13g2_decap_8
XFILLER_40_1019 VDD VSS sg13g2_decap_8
XFILLER_57_323 VDD VSS sg13g2_decap_8
XFILLER_100_987 VDD VSS sg13g2_decap_8
XFILLER_84_142 VDD VSS sg13g2_decap_8
XFILLER_27_35 VDD VSS sg13g2_decap_8
XFILLER_45_518 VDD VSS sg13g2_decap_8
XFILLER_100_998 VDD VSS sg13g2_fill_1
XFILLER_26_721 VDD VSS sg13g2_decap_8
XFILLER_72_359 VDD VSS sg13g2_decap_8
XFILLER_25_231 VDD VSS sg13g2_decap_8
XFILLER_81_893 VDD VSS sg13g2_decap_8
XFILLER_53_573 VDD VSS sg13g2_decap_8
XFILLER_41_713 VDD VSS sg13g2_decap_8
XFILLER_26_798 VDD VSS sg13g2_decap_8
XFILLER_14_938 VDD VSS sg13g2_decap_8
XFILLER_13_448 VDD VSS sg13g2_decap_8
XFILLER_43_56 VDD VSS sg13g2_decap_8
XFILLER_5_658 VDD VSS sg13g2_decap_8
XFILLER_107_597 VDD VSS sg13g2_decap_8
XFILLER_4_168 VDD VSS sg13g2_decap_8
XFILLER_4_28 VDD VSS sg13g2_decap_8
XFILLER_68_42 VDD VSS sg13g2_decap_8
XFILLER_110_718 VDD VSS sg13g2_decap_8
XFILLER_103_770 VDD VSS sg13g2_decap_8
XFILLER_76_610 VDD VSS sg13g2_decap_8
XFILLER_1_875 VDD VSS sg13g2_decap_8
XFILLER_68_75 VDD VSS sg13g2_decap_8
XFILLER_76_632 VDD VSS sg13g2_decap_8
XFILLER_76_643 VDD VSS sg13g2_decap_8
XFILLER_76_621 VDD VSS sg13g2_fill_1
XFILLER_88_492 VDD VSS sg13g2_decap_4
XFILLER_0_385 VDD VSS sg13g2_decap_8
XFILLER_64_816 VDD VSS sg13g2_decap_8
XFILLER_63_304 VDD VSS sg13g2_decap_8
XFILLER_36_518 VDD VSS sg13g2_decap_8
XFILLER_48_367 VDD VSS sg13g2_decap_8
X_2304__95 VDD VSS _2304__95/L_HI sg13g2_tiehi
XFILLER_90_112 VDD VSS sg13g2_decap_8
XFILLER_84_63 VDD VSS sg13g2_decap_8
XFILLER_29_581 VDD VSS sg13g2_decap_8
XFILLER_17_721 VDD VSS sg13g2_decap_8
XFILLER_63_359 VDD VSS sg13g2_decap_8
XFILLER_16_231 VDD VSS sg13g2_decap_8
XFILLER_1_1057 VDD VSS sg13g2_decap_4
XFILLER_90_167 VDD VSS sg13g2_decap_8
XFILLER_17_798 VDD VSS sg13g2_decap_8
XFILLER_90_7 VDD VSS sg13g2_decap_8
XFILLER_32_735 VDD VSS sg13g2_decap_8
XFILLER_31_245 VDD VSS sg13g2_decap_8
XFILLER_9_931 VDD VSS sg13g2_decap_8
X_1701_ _1725_/A _1701_/B _1701_/Y VDD VSS sg13g2_nor2_1
XFILLER_8_441 VDD VSS sg13g2_decap_8
X_1632_ _1639_/A _1632_/B _1632_/Y VDD VSS sg13g2_nor2_1
X_1563_ _1577_/S0 _2240_/Q _2232_/Q _2224_/Q _2216_/Q _2287_/Q _1564_/A VDD VSS sg13g2_mux4_1
X_1494_ _2101_/A _1494_/B _2266_/D VDD VSS sg13g2_nor2_1
XFILLER_98_267 VDD VSS sg13g2_decap_8
XFILLER_95_952 VDD VSS sg13g2_decap_8
XFILLER_67_621 VDD VSS sg13g2_decap_8
XFILLER_94_440 VDD VSS sg13g2_decap_8
XFILLER_12_0 VDD VSS sg13g2_decap_8
XFILLER_66_153 VDD VSS sg13g2_decap_8
XFILLER_27_518 VDD VSS sg13g2_decap_8
XFILLER_39_345 VDD VSS sg13g2_decap_8
XFILLER_82_646 VDD VSS sg13g2_decap_8
X_2115_ _2115_/A _2115_/B _2366_/D VDD VSS sg13g2_nor2_1
XFILLER_67_698 VDD VSS sg13g2_decap_8
XFILLER_70_808 VDD VSS sg13g2_decap_8
X_2046_ _2156_/A _2040_/A _2329_/D VDD VSS sg13g2_nor2b_1
XFILLER_54_359 VDD VSS sg13g2_decap_8
XFILLER_54_348 VDD VSS sg13g2_decap_4
XFILLER_63_860 VDD VSS sg13g2_decap_8
Xfanout38 _1338_/A2 _1322_/A2 VDD VSS sg13g2_buf_1
Xfanout16 _1342_/B1 _1482_/B1 VDD VSS sg13g2_buf_1
XFILLER_35_595 VDD VSS sg13g2_decap_8
XFILLER_23_735 VDD VSS sg13g2_decap_8
Xfanout27 _1448_/X _1453_/B VDD VSS sg13g2_buf_1
XFILLER_50_532 VDD VSS sg13g2_decap_8
Xfanout49 _2308_/Q _1724_/S VDD VSS sg13g2_buf_1
XFILLER_22_245 VDD VSS sg13g2_decap_8
Xhold452 _2239_/Q VDD VSS hold452/X sg13g2_dlygate4sd3_1
X_2164__212 VDD VSS _2164_/RESET_B sg13g2_tiehi
Xhold430 _1648_/Y VDD VSS _1649_/B sg13g2_dlygate4sd3_1
Xhold441 _2364_/Q VDD VSS _1501_/B sg13g2_dlygate4sd3_1
XFILLER_1_105 VDD VSS sg13g2_decap_8
Xhold463 _2280_/Q VDD VSS hold463/X sg13g2_dlygate4sd3_1
Xhold474 _1722_/Y VDD VSS _2319_/D sg13g2_dlygate4sd3_1
XFILLER_104_545 VDD VSS sg13g2_fill_1
XFILLER_104_556 VDD VSS sg13g2_decap_8
Xhold496 _2352_/Q VDD VSS _2099_/A sg13g2_dlygate4sd3_1
Xhold485 _1575_/Y VDD VSS _1576_/B sg13g2_dlygate4sd3_1
XFILLER_86_930 VDD VSS sg13g2_decap_8
XFILLER_85_440 VDD VSS sg13g2_decap_8
XFILLER_58_665 VDD VSS sg13g2_decap_8
XFILLER_38_56 VDD VSS sg13g2_decap_8
XFILLER_86_996 VDD VSS sg13g2_decap_8
XFILLER_46_838 VDD VSS sg13g2_fill_2
XFILLER_57_186 VDD VSS sg13g2_decap_8
XFILLER_18_518 VDD VSS sg13g2_decap_8
XFILLER_45_315 VDD VSS sg13g2_decap_8
XFILLER_79_1059 VDD VSS sg13g2_fill_2
XFILLER_73_646 VDD VSS sg13g2_decap_8
XFILLER_72_189 VDD VSS sg13g2_decap_8
XFILLER_54_871 VDD VSS sg13g2_decap_8
XFILLER_41_543 VDD VSS sg13g2_decap_8
XFILLER_26_595 VDD VSS sg13g2_decap_8
XFILLER_14_735 VDD VSS sg13g2_decap_8
XFILLER_54_99 VDD VSS sg13g2_decap_8
XFILLER_13_245 VDD VSS sg13g2_decap_8
XFILLER_70_21 VDD VSS sg13g2_decap_8
XFILLER_41_587 VDD VSS sg13g2_decap_8
XFILLER_9_238 VDD VSS sg13g2_decap_8
XFILLER_16_1043 VDD VSS sg13g2_decap_8
XFILLER_10_952 VDD VSS sg13g2_decap_8
XFILLER_103_1057 VDD VSS sg13g2_decap_4
XFILLER_70_98 VDD VSS sg13g2_decap_8
XFILLER_6_945 VDD VSS sg13g2_decap_8
XFILLER_5_455 VDD VSS sg13g2_decap_8
XFILLER_79_63 VDD VSS sg13g2_decap_8
XFILLER_110_515 VDD VSS sg13g2_decap_8
XFILLER_95_248 VDD VSS sg13g2_decap_8
XFILLER_62_1052 VDD VSS sg13g2_decap_8
XFILLER_1_672 VDD VSS sg13g2_decap_8
XFILLER_76_462 VDD VSS sg13g2_decap_8
XFILLER_95_84 VDD VSS sg13g2_decap_8
XFILLER_23_1036 VDD VSS sg13g2_decap_8
XFILLER_37_805 VDD VSS sg13g2_decap_8
XFILLER_0_182 VDD VSS sg13g2_decap_8
XFILLER_92_922 VDD VSS sg13g2_fill_1
XFILLER_91_410 VDD VSS sg13g2_decap_4
XFILLER_64_613 VDD VSS sg13g2_decap_8
XFILLER_36_315 VDD VSS sg13g2_decap_8
XFILLER_48_175 VDD VSS sg13g2_decap_8
XFILLER_91_454 VDD VSS sg13g2_decap_8
XFILLER_63_145 VDD VSS sg13g2_decap_8
XFILLER_45_882 VDD VSS sg13g2_decap_8
XFILLER_91_498 VDD VSS sg13g2_fill_1
XFILLER_17_595 VDD VSS sg13g2_decap_8
XFILLER_32_532 VDD VSS sg13g2_decap_8
XFILLER_44_392 VDD VSS sg13g2_decap_8
XFILLER_20_749 VDD VSS sg13g2_decap_8
XFILLER_30_1029 VDD VSS sg13g2_decap_8
XFILLER_105_309 VDD VSS sg13g2_decap_8
X_1615_ _1639_/A _1615_/B _1615_/Y VDD VSS sg13g2_nor2_1
X_1546_ _1545_/Y VDD _1546_/Y VSS _1592_/A _1543_/Y sg13g2_o21ai_1
XFILLER_99_576 VDD VSS sg13g2_decap_8
XFILLER_87_738 VDD VSS sg13g2_decap_8
XFILLER_8_1008 VDD VSS sg13g2_decap_8
XFILLER_101_548 VDD VSS sg13g2_fill_2
XFILLER_86_237 VDD VSS sg13g2_decap_8
X_1477_ VSS VDD _1196_/Y _1479_/A2 _2257_/D _1476_/Y sg13g2_a21oi_1
XFILLER_28_805 VDD VSS sg13g2_decap_8
XFILLER_55_613 VDD VSS sg13g2_decap_8
XFILLER_27_315 VDD VSS sg13g2_decap_8
XFILLER_39_175 VDD VSS sg13g2_decap_8
XFILLER_82_443 VDD VSS sg13g2_decap_8
XFILLER_82_454 VDD VSS sg13g2_fill_2
XFILLER_54_134 VDD VSS sg13g2_decap_8
XFILLER_70_605 VDD VSS sg13g2_decap_8
XFILLER_36_882 VDD VSS sg13g2_decap_8
XFILLER_42_318 VDD VSS sg13g2_decap_8
X_2029_ _2021_/X _2040_/A _2036_/S _2030_/B VDD VSS sg13g2_mux2_1
XFILLER_39_1032 VDD VSS sg13g2_decap_8
XFILLER_54_189 VDD VSS sg13g2_decap_8
XFILLER_24_14 VDD VSS sg13g2_decap_8
XFILLER_23_532 VDD VSS sg13g2_decap_8
XFILLER_35_392 VDD VSS sg13g2_decap_8
XFILLER_51_874 VDD VSS sg13g2_decap_4
XFILLER_11_749 VDD VSS sg13g2_decap_8
XFILLER_10_259 VDD VSS sg13g2_decap_8
XFILLER_50_395 VDD VSS sg13g2_decap_8
XFILLER_109_637 VDD VSS sg13g2_decap_8
XFILLER_40_35 VDD VSS sg13g2_decap_8
XFILLER_108_147 VDD VSS sg13g2_decap_8
XFILLER_105_854 VDD VSS sg13g2_decap_8
XFILLER_46_1003 VDD VSS sg13g2_decap_8
XFILLER_3_959 VDD VSS sg13g2_decap_8
XFILLER_104_342 VDD VSS sg13g2_decap_8
Xhold293 _2362_/Q VDD VSS _1500_/D sg13g2_dlygate4sd3_1
XFILLER_2_469 VDD VSS sg13g2_decap_8
XFILLER_86_760 VDD VSS sg13g2_decap_8
XFILLER_19_805 VDD VSS sg13g2_decap_8
XFILLER_74_933 VDD VSS sg13g2_decap_8
XFILLER_100_581 VDD VSS sg13g2_decap_8
XFILLER_59_985 VDD VSS sg13g2_decap_8
XFILLER_18_315 VDD VSS sg13g2_decap_8
XFILLER_65_21 VDD VSS sg13g2_decap_8
XFILLER_85_292 VDD VSS sg13g2_decap_8
XFILLER_73_421 VDD VSS sg13g2_decap_8
XFILLER_45_112 VDD VSS sg13g2_decap_4
XFILLER_34_819 VDD VSS sg13g2_decap_8
XFILLER_27_882 VDD VSS sg13g2_decap_8
XFILLER_65_87 VDD VSS sg13g2_decap_8
XFILLER_92_1023 VDD VSS sg13g2_fill_2
XFILLER_92_1012 VDD VSS sg13g2_decap_8
XFILLER_73_498 VDD VSS sg13g2_decap_8
XFILLER_14_532 VDD VSS sg13g2_decap_8
XFILLER_26_392 VDD VSS sg13g2_decap_8
XFILLER_33_329 VDD VSS sg13g2_decap_8
XFILLER_45_189 VDD VSS sg13g2_decap_8
XFILLER_92_1056 VDD VSS sg13g2_decap_4
XFILLER_81_42 VDD VSS sg13g2_decap_8
XFILLER_53_1018 VDD VSS sg13g2_fill_2
XFILLER_42_896 VDD VSS sg13g2_decap_8
XFILLER_41_395 VDD VSS sg13g2_decap_8
XFILLER_14_91 VDD VSS sg13g2_decap_8
XFILLER_6_742 VDD VSS sg13g2_decap_8
XFILLER_5_252 VDD VSS sg13g2_decap_8
XFILLER_53_7 VDD VSS sg13g2_decap_8
X_1400_ VDD _2222_/D _1400_/A VSS sg13g2_inv_1
XFILLER_69_727 VDD VSS sg13g2_decap_8
XFILLER_68_204 VDD VSS sg13g2_decap_8
XFILLER_110_301 VDD VSS sg13g2_decap_8
XFILLER_96_535 VDD VSS sg13g2_decap_4
X_1331_ VDD _2195_/D _1331_/A VSS sg13g2_inv_1
XFILLER_111_868 VDD VSS sg13g2_decap_8
XFILLER_96_557 VDD VSS sg13g2_decap_8
XFILLER_77_760 VDD VSS sg13g2_decap_8
X_1262_ _1234_/B _1236_/C _1235_/A _1262_/X VDD VSS sg13g2_a21o_1
XFILLER_49_440 VDD VSS sg13g2_decap_8
XFILLER_110_389 VDD VSS sg13g2_decap_8
XFILLER_37_602 VDD VSS sg13g2_decap_8
XFILLER_65_944 VDD VSS sg13g2_decap_8
X_1193_ VDD _1193_/Y _1487_/A VSS sg13g2_inv_1
XFILLER_36_112 VDD VSS sg13g2_decap_8
X_2293__137 VDD VSS _2293_/RESET_B sg13g2_tiehi
X_2258__235 VDD VSS _2258_/RESET_B sg13g2_tiehi
XFILLER_92_763 VDD VSS sg13g2_decap_8
XFILLER_91_262 VDD VSS sg13g2_decap_8
XFILLER_37_679 VDD VSS sg13g2_decap_8
XFILLER_25_819 VDD VSS sg13g2_decap_8
XFILLER_64_465 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_52_638 VDD VSS sg13g2_decap_8
XFILLER_45_690 VDD VSS sg13g2_decap_8
XFILLER_18_882 VDD VSS sg13g2_decap_8
XFILLER_51_126 VDD VSS sg13g2_decap_8
XFILLER_24_329 VDD VSS sg13g2_decap_8
XFILLER_36_189 VDD VSS sg13g2_decap_8
XFILLER_17_392 VDD VSS sg13g2_decap_8
XFILLER_60_682 VDD VSS sg13g2_decap_4
XFILLER_33_896 VDD VSS sg13g2_decap_8
XFILLER_20_546 VDD VSS sg13g2_decap_8
XFILLER_106_629 VDD VSS sg13g2_decap_8
Xin_data_pads\[0\].in_data_pad IOVDD IOVSS _1364_/A in_data_PADs[0] VDD VSS sg13g2_IOPadIn
XFILLER_10_49 VDD VSS sg13g2_decap_8
XFILLER_102_802 VDD VSS sg13g2_decap_4
XFILLER_102_846 VDD VSS sg13g2_decap_8
XFILLER_101_323 VDD VSS sg13g2_decap_8
XFILLER_99_373 VDD VSS sg13g2_decap_8
X_1529_ VDD _1529_/Y _1529_/A VSS sg13g2_inv_1
XFILLER_59_215 VDD VSS sg13g2_decap_8
XFILLER_19_14 VDD VSS sg13g2_decap_8
XFILLER_68_771 VDD VSS sg13g2_decap_8
XFILLER_28_602 VDD VSS sg13g2_decap_8
XFILLER_27_112 VDD VSS sg13g2_decap_8
XFILLER_71_914 VDD VSS sg13g2_decap_8
XFILLER_56_977 VDD VSS sg13g2_decap_8
XFILLER_28_679 VDD VSS sg13g2_decap_8
XFILLER_16_819 VDD VSS sg13g2_decap_8
XFILLER_70_435 VDD VSS sg13g2_decap_8
XFILLER_55_487 VDD VSS sg13g2_decap_8
XFILLER_15_329 VDD VSS sg13g2_decap_8
XFILLER_35_35 VDD VSS sg13g2_decap_8
XFILLER_42_126 VDD VSS sg13g2_decap_8
XFILLER_27_189 VDD VSS sg13g2_decap_8
XFILLER_51_682 VDD VSS sg13g2_decap_8
XFILLER_24_896 VDD VSS sg13g2_decap_8
XFILLER_11_546 VDD VSS sg13g2_decap_8
XFILLER_51_23 VDD VSS sg13g2_fill_1
XFILLER_50_181 VDD VSS sg13g2_decap_8
XFILLER_7_539 VDD VSS sg13g2_decap_8
XFILLER_51_67 VDD VSS sg13g2_decap_8
XFILLER_109_434 VDD VSS sg13g2_decap_8
XFILLER_13_1057 VDD VSS sg13g2_decap_4
XFILLER_105_651 VDD VSS sg13g2_decap_8
XFILLER_3_756 VDD VSS sg13g2_decap_8
XFILLER_2_266 VDD VSS sg13g2_decap_8
XFILLER_93_505 VDD VSS sg13g2_decap_8
XFILLER_76_42 VDD VSS sg13g2_decap_8
XFILLER_47_922 VDD VSS sg13g2_decap_8
XFILLER_59_782 VDD VSS sg13g2_decap_8
XFILLER_19_602 VDD VSS sg13g2_decap_8
XFILLER_101_890 VDD VSS sg13g2_fill_1
XFILLER_58_281 VDD VSS sg13g2_decap_8
XFILLER_18_112 VDD VSS sg13g2_decap_8
XFILLER_47_999 VDD VSS sg13g2_decap_8
XFILLER_34_616 VDD VSS sg13g2_decap_8
XFILLER_19_679 VDD VSS sg13g2_decap_8
XFILLER_92_63 VDD VSS sg13g2_decap_8
XFILLER_18_189 VDD VSS sg13g2_decap_8
XFILLER_33_126 VDD VSS sg13g2_decap_8
XFILLER_61_446 VDD VSS sg13g2_decap_8
XFILLER_15_896 VDD VSS sg13g2_decap_8
X_1880_ _1880_/Y _1880_/A _1880_/B VDD VSS sg13g2_xnor2_1
XFILLER_42_693 VDD VSS sg13g2_decap_8
XFILLER_30_833 VDD VSS sg13g2_decap_8
XFILLER_41_181 VDD VSS sg13g2_decap_8
X_2363_ _2363_/RESET_B VSS VDD _2363_/D _2363_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_111_665 VDD VSS sg13g2_decap_8
XFILLER_97_888 VDD VSS sg13g2_decap_8
XFILLER_69_579 VDD VSS sg13g2_decap_8
XFILLER_96_343 VDD VSS sg13g2_decap_8
X_1314_ _1314_/Y _1482_/B1 hold338/X _1482_/A2 _2374_/Q VDD VSS sg13g2_a22oi_1
XFILLER_99_1018 VDD VSS sg13g2_fill_1
XFILLER_99_1007 VDD VSS sg13g2_decap_8
XFILLER_110_175 VDD VSS sg13g2_decap_8
XFILLER_38_933 VDD VSS sg13g2_decap_8
X_2294_ _2294_/RESET_B VSS VDD _2294_/D _2294_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_65_752 VDD VSS sg13g2_decap_8
X_1245_ _1247_/D _2291_/Q _2253_/Q VDD VSS sg13g2_xnor2_1
XFILLER_49_281 VDD VSS sg13g2_decap_8
XFILLER_53_925 VDD VSS sg13g2_decap_4
XFILLER_25_616 VDD VSS sg13g2_decap_8
XFILLER_64_240 VDD VSS sg13g2_decap_8
XFILLER_37_476 VDD VSS sg13g2_decap_8
XFILLER_52_424 VDD VSS sg13g2_decap_8
XFILLER_24_126 VDD VSS sg13g2_decap_8
XFILLER_53_969 VDD VSS sg13g2_decap_8
XFILLER_80_788 VDD VSS sg13g2_fill_1
XFILLER_36_1057 VDD VSS sg13g2_decap_4
XFILLER_33_693 VDD VSS sg13g2_decap_8
XFILLER_21_833 VDD VSS sg13g2_decap_8
XFILLER_20_343 VDD VSS sg13g2_decap_8
XFILLER_107_905 VDD VSS sg13g2_decap_8
XFILLER_82_1033 VDD VSS sg13g2_decap_8
XFILLER_88_844 VDD VSS sg13g2_decap_8
XFILLER_99_170 VDD VSS sg13g2_decap_8
XFILLER_43_1017 VDD VSS sg13g2_decap_8
XFILLER_48_708 VDD VSS sg13g2_decap_8
XFILLER_75_549 VDD VSS sg13g2_fill_1
XFILLER_29_966 VDD VSS sg13g2_decap_8
XFILLER_56_763 VDD VSS sg13g2_decap_8
XFILLER_44_914 VDD VSS sg13g2_decap_8
XFILLER_16_616 VDD VSS sg13g2_decap_8
XFILLER_46_56 VDD VSS sg13g2_decap_8
XFILLER_28_476 VDD VSS sg13g2_decap_8
XFILLER_83_571 VDD VSS sg13g2_decap_8
XFILLER_55_273 VDD VSS sg13g2_decap_8
XFILLER_15_126 VDD VSS sg13g2_decap_8
XFILLER_43_413 VDD VSS sg13g2_decap_8
XFILLER_71_777 VDD VSS sg13g2_decap_8
XFILLER_71_755 VDD VSS sg13g2_fill_2
XFILLER_102_84 VDD VSS sg13g2_decap_8
XFILLER_24_693 VDD VSS sg13g2_decap_8
XFILLER_51_490 VDD VSS sg13g2_decap_4
XFILLER_12_833 VDD VSS sg13g2_decap_8
XFILLER_62_77 VDD VSS sg13g2_decap_8
X_2172__196 VDD VSS _2172_/RESET_B sg13g2_tiehi
XFILLER_11_343 VDD VSS sg13g2_decap_8
XFILLER_7_28 VDD VSS sg13g2_decap_8
XFILLER_8_826 VDD VSS sg13g2_decap_8
XFILLER_7_336 VDD VSS sg13g2_decap_8
XFILLER_109_286 VDD VSS sg13g2_fill_2
XFILLER_98_619 VDD VSS sg13g2_decap_8
XFILLER_11_70 VDD VSS sg13g2_decap_8
XFILLER_3_553 VDD VSS sg13g2_decap_8
XFILLER_106_993 VDD VSS sg13g2_decap_8
XFILLER_79_844 VDD VSS sg13g2_fill_1
XFILLER_105_470 VDD VSS sg13g2_fill_1
XFILLER_87_63 VDD VSS sg13g2_decap_8
XFILLER_94_836 VDD VSS sg13g2_decap_8
XFILLER_79_888 VDD VSS sg13g2_decap_8
XFILLER_66_505 VDD VSS sg13g2_decap_8
XFILLER_93_324 VDD VSS sg13g2_fill_2
XFILLER_47_730 VDD VSS sg13g2_fill_2
XFILLER_16_7 VDD VSS sg13g2_decap_8
XFILLER_4_1022 VDD VSS sg13g2_decap_8
XFILLER_74_560 VDD VSS sg13g2_decap_8
XFILLER_59_1013 VDD VSS sg13g2_decap_8
XFILLER_62_700 VDD VSS sg13g2_fill_2
XFILLER_35_903 VDD VSS sg13g2_decap_8
XFILLER_59_1024 VDD VSS sg13g2_decap_4
XFILLER_62_733 VDD VSS sg13g2_decap_8
XFILLER_19_476 VDD VSS sg13g2_decap_8
XFILLER_34_413 VDD VSS sg13g2_decap_8
XFILLER_46_284 VDD VSS sg13g2_decap_8
XFILLER_50_939 VDD VSS sg13g2_decap_8
XFILLER_61_287 VDD VSS sg13g2_decap_8
X_1932_ _1933_/A _1933_/B _1932_/Y VDD VSS sg13g2_nor2b_1
XFILLER_30_630 VDD VSS sg13g2_decap_8
XFILLER_15_693 VDD VSS sg13g2_decap_8
X_1863_ _1892_/B _1863_/A _1863_/B VDD VSS sg13g2_xnor2_1
X_1794_ _1801_/B _2224_/Q _2216_/Q VDD VSS sg13g2_nand2b_1
XFILLER_104_908 VDD VSS sg13g2_decap_8
XFILLER_66_1028 VDD VSS sg13g2_decap_8
XFILLER_42_0 VDD VSS sg13g2_decap_8
XFILLER_112_952 VDD VSS sg13g2_decap_8
X_2346_ _2346_/RESET_B VSS VDD _2346_/D _2346_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_111_462 VDD VSS sg13g2_decap_8
XFILLER_84_313 VDD VSS sg13g2_decap_4
XFILLER_96_140 VDD VSS sg13g2_decap_8
XFILLER_42_1050 VDD VSS sg13g2_decap_8
XFILLER_38_730 VDD VSS sg13g2_decap_8
X_2277_ _2277_/RESET_B VSS VDD _2277_/D _2277_/Q clkload0/A sg13g2_dfrbpq_1
X_1228_ _1228_/A _1228_/B _2365_/D VDD VSS sg13g2_nor2_1
XFILLER_26_903 VDD VSS sg13g2_decap_8
XFILLER_93_880 VDD VSS sg13g2_decap_4
XFILLER_53_711 VDD VSS sg13g2_decap_8
XFILLER_25_413 VDD VSS sg13g2_decap_8
XFILLER_37_273 VDD VSS sg13g2_decap_8
XFILLER_80_530 VDD VSS sg13g2_decap_8
XFILLER_52_243 VDD VSS sg13g2_decap_8
XFILLER_34_980 VDD VSS sg13g2_decap_8
XFILLER_40_405 VDD VSS sg13g2_decap_8
XFILLER_21_630 VDD VSS sg13g2_decap_8
XFILLER_33_490 VDD VSS sg13g2_decap_8
XFILLER_20_140 VDD VSS sg13g2_decap_8
XFILLER_32_14 VDD VSS sg13g2_decap_8
XFILLER_107_702 VDD VSS sg13g2_decap_8
XFILLER_107_779 VDD VSS sg13g2_decap_8
XFILLER_106_245 VDD VSS sg13g2_decap_8
XFILLER_103_952 VDD VSS sg13g2_decap_8
XFILLER_87_151 VDD VSS sg13g2_decap_8
XFILLER_0_567 VDD VSS sg13g2_decap_8
XFILLER_76_858 VDD VSS sg13g2_decap_8
XFILLER_102_484 VDD VSS sg13g2_decap_8
XFILLER_75_313 VDD VSS sg13g2_decap_8
XFILLER_90_305 VDD VSS sg13g2_decap_8
XFILLER_29_763 VDD VSS sg13g2_decap_8
XFILLER_17_903 VDD VSS sg13g2_decap_8
XFILLER_57_99 VDD VSS sg13g2_fill_1
XFILLER_57_88 VDD VSS sg13g2_decap_8
XFILLER_73_21 VDD VSS sg13g2_decap_8
XFILLER_56_560 VDD VSS sg13g2_decap_8
XFILLER_44_711 VDD VSS sg13g2_decap_8
XFILLER_16_413 VDD VSS sg13g2_decap_8
XFILLER_28_273 VDD VSS sg13g2_decap_8
XFILLER_43_210 VDD VSS sg13g2_decap_8
XFILLER_73_98 VDD VSS sg13g2_decap_8
XFILLER_32_917 VDD VSS sg13g2_decap_8
XFILLER_25_980 VDD VSS sg13g2_decap_8
XFILLER_44_788 VDD VSS sg13g2_decap_8
XFILLER_44_799 VDD VSS sg13g2_fill_1
XFILLER_43_265 VDD VSS sg13g2_decap_8
XFILLER_106_1000 VDD VSS sg13g2_decap_8
XFILLER_12_630 VDD VSS sg13g2_decap_8
XFILLER_24_490 VDD VSS sg13g2_decap_8
XFILLER_31_427 VDD VSS sg13g2_decap_8
XFILLER_11_140 VDD VSS sg13g2_decap_8
XFILLER_89_1017 VDD VSS sg13g2_decap_8
XFILLER_8_623 VDD VSS sg13g2_decap_8
XFILLER_7_133 VDD VSS sg13g2_decap_8
XFILLER_22_91 VDD VSS sg13g2_decap_8
XFILLER_4_840 VDD VSS sg13g2_decap_8
XFILLER_98_84 VDD VSS sg13g2_decap_8
XFILLER_3_350 VDD VSS sg13g2_decap_8
XFILLER_106_790 VDD VSS sg13g2_decap_8
X_2200_ _2200_/RESET_B VSS VDD _2200_/D _2200_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_112_259 VDD VSS sg13g2_decap_8
XFILLER_65_1050 VDD VSS sg13g2_decap_8
XFILLER_26_1001 VDD VSS sg13g2_decap_8
XFILLER_79_685 VDD VSS sg13g2_decap_8
XFILLER_78_140 VDD VSS sg13g2_decap_8
X_2131_ _2131_/A _2131_/B _2369_/D VDD VSS sg13g2_nor2_1
XFILLER_94_622 VDD VSS sg13g2_decap_8
XFILLER_67_858 VDD VSS sg13g2_fill_2
XFILLER_39_549 VDD VSS sg13g2_decap_8
XFILLER_94_655 VDD VSS sg13g2_decap_8
XFILLER_82_806 VDD VSS sg13g2_decap_8
X_2062_ _2066_/A _2062_/B _2025_/A VDD VSS sg13g2_nand2b_1
XFILLER_81_305 VDD VSS sg13g2_decap_8
XFILLER_93_154 VDD VSS sg13g2_decap_8
XFILLER_94_699 VDD VSS sg13g2_decap_8
XFILLER_93_198 VDD VSS sg13g2_decap_8
XFILLER_93_165 VDD VSS sg13g2_fill_2
XFILLER_47_571 VDD VSS sg13g2_fill_1
XFILLER_35_700 VDD VSS sg13g2_decap_8
XFILLER_19_273 VDD VSS sg13g2_decap_8
XFILLER_34_210 VDD VSS sg13g2_decap_8
XFILLER_90_872 VDD VSS sg13g2_fill_2
XFILLER_23_917 VDD VSS sg13g2_decap_8
XFILLER_50_703 VDD VSS sg13g2_fill_2
XFILLER_50_725 VDD VSS sg13g2_fill_2
XFILLER_35_777 VDD VSS sg13g2_decap_8
XFILLER_16_980 VDD VSS sg13g2_decap_8
XFILLER_72_1032 VDD VSS sg13g2_decap_8
XFILLER_15_490 VDD VSS sg13g2_decap_8
XFILLER_22_427 VDD VSS sg13g2_decap_8
XFILLER_34_287 VDD VSS sg13g2_decap_8
X_1915_ _1917_/A _1915_/A _1915_/B VDD VSS sg13g2_xnor2_1
Xclkbuf_leaf_14_clk clkbuf_2_2__f_clk/X _2373_/CLK VDD VSS sg13g2_buf_8
XFILLER_31_994 VDD VSS sg13g2_decap_8
X_1846_ VDD _1846_/Y _1856_/A VSS sg13g2_inv_1
X_1777_ _1777_/Y _2214_/Q _2222_/Q VDD VSS sg13g2_nand2b_1
XFILLER_89_405 VDD VSS sg13g2_decap_8
XFILLER_98_983 VDD VSS sg13g2_decap_8
XFILLER_100_911 VDD VSS sg13g2_decap_8
XFILLER_69_195 VDD VSS sg13g2_decap_4
XFILLER_69_184 VDD VSS sg13g2_decap_8
X_2329_ _2329_/RESET_B VSS VDD _2329_/D _2329_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_100_966 VDD VSS sg13g2_decap_8
XFILLER_58_869 VDD VSS sg13g2_fill_2
XFILLER_27_14 VDD VSS sg13g2_decap_8
XFILLER_73_839 VDD VSS sg13g2_decap_8
XFILLER_72_338 VDD VSS sg13g2_decap_8
XFILLER_26_700 VDD VSS sg13g2_decap_8
XFILLER_84_198 VDD VSS sg13g2_decap_4
XFILLER_25_210 VDD VSS sg13g2_decap_8
X_2238__266 VDD VSS _2238_/RESET_B sg13g2_tiehi
XFILLER_26_777 VDD VSS sg13g2_decap_8
XFILLER_14_917 VDD VSS sg13g2_decap_8
XFILLER_13_427 VDD VSS sg13g2_decap_8
XFILLER_43_35 VDD VSS sg13g2_decap_8
XFILLER_25_287 VDD VSS sg13g2_decap_8
XFILLER_40_224 VDD VSS sg13g2_fill_1
XFILLER_41_769 VDD VSS sg13g2_decap_8
XFILLER_22_994 VDD VSS sg13g2_decap_8
XFILLER_5_637 VDD VSS sg13g2_decap_8
XFILLER_4_147 VDD VSS sg13g2_decap_8
XFILLER_107_576 VDD VSS sg13g2_decap_8
XFILLER_49_1056 VDD VSS sg13g2_decap_4
XFILLER_89_950 VDD VSS sg13g2_decap_8
XFILLER_1_854 VDD VSS sg13g2_decap_8
XFILLER_68_21 VDD VSS sg13g2_decap_8
XFILLER_89_972 VDD VSS sg13g2_decap_8
XFILLER_49_825 VDD VSS sg13g2_decap_8
XFILLER_0_364 VDD VSS sg13g2_decap_8
XFILLER_68_65 VDD VSS sg13g2_fill_1
XFILLER_48_302 VDD VSS sg13g2_decap_8
XFILLER_88_471 VDD VSS sg13g2_decap_8
XFILLER_75_154 VDD VSS sg13g2_decap_8
XFILLER_48_357 VDD VSS sg13g2_fill_2
XFILLER_76_699 VDD VSS sg13g2_decap_8
XFILLER_84_42 VDD VSS sg13g2_decap_8
XFILLER_75_165 VDD VSS sg13g2_fill_2
XFILLER_57_880 VDD VSS sg13g2_decap_8
XFILLER_29_560 VDD VSS sg13g2_decap_8
XFILLER_17_700 VDD VSS sg13g2_decap_8
XFILLER_95_1043 VDD VSS sg13g2_decap_8
XFILLER_91_658 VDD VSS sg13g2_decap_4
XFILLER_91_669 VDD VSS sg13g2_decap_8
XFILLER_90_146 VDD VSS sg13g2_decap_8
XFILLER_63_338 VDD VSS sg13g2_decap_8
XFILLER_16_210 VDD VSS sg13g2_decap_8
XFILLER_1_1036 VDD VSS sg13g2_decap_8
XFILLER_32_714 VDD VSS sg13g2_decap_8
XFILLER_17_91 VDD VSS sg13g2_decap_8
XFILLER_17_777 VDD VSS sg13g2_decap_8
XFILLER_71_371 VDD VSS sg13g2_decap_8
XFILLER_44_585 VDD VSS sg13g2_decap_8
XFILLER_16_287 VDD VSS sg13g2_decap_8
XFILLER_31_224 VDD VSS sg13g2_decap_8
XFILLER_9_910 VDD VSS sg13g2_decap_8
XFILLER_83_7 VDD VSS sg13g2_decap_8
XFILLER_8_420 VDD VSS sg13g2_decap_8
XFILLER_13_994 VDD VSS sg13g2_decap_8
X_2289__153 VDD VSS _2289_/RESET_B sg13g2_tiehi
X_1700_ _1699_/Y VDD _1700_/Y VSS _1720_/A hold466/X sg13g2_o21ai_1
XFILLER_9_987 VDD VSS sg13g2_decap_8
XFILLER_8_497 VDD VSS sg13g2_decap_8
X_1631_ _1630_/Y VDD _1631_/Y VSS _1634_/A hold532/X sg13g2_o21ai_1
XFILLER_99_736 VDD VSS sg13g2_fill_2
X_1562_ _1576_/A _1562_/B _2279_/D VDD VSS sg13g2_nor2_1
XFILLER_98_246 VDD VSS sg13g2_decap_8
X_1493_ _1493_/A _1493_/B _1494_/B VDD VSS sg13g2_nor2_1
XFILLER_86_419 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_3_clk clkbuf_leaf_5_clk/A _2245_/CLK VDD VSS sg13g2_buf_8
XFILLER_95_931 VDD VSS sg13g2_decap_8
XFILLER_79_493 VDD VSS sg13g2_fill_2
XFILLER_79_482 VDD VSS sg13g2_decap_8
XFILLER_39_324 VDD VSS sg13g2_decap_8
X_2114_ _1688_/B VDD _2115_/B VSS _1259_/A hold566/X sg13g2_o21ai_1
XFILLER_67_677 VDD VSS sg13g2_decap_8
XFILLER_82_625 VDD VSS sg13g2_decap_8
XFILLER_94_496 VDD VSS sg13g2_decap_8
XFILLER_55_839 VDD VSS sg13g2_decap_8
XFILLER_48_891 VDD VSS sg13g2_decap_4
XFILLER_54_327 VDD VSS sg13g2_decap_8
X_2045_ VDD _2328_/D _2045_/A VSS sg13g2_inv_1
XFILLER_81_157 VDD VSS sg13g2_decap_8
XFILLER_35_574 VDD VSS sg13g2_decap_8
XFILLER_23_714 VDD VSS sg13g2_decap_8
Xfanout28 _1428_/Y _1429_/B VDD VSS sg13g2_buf_1
Xfanout17 fanout22/X _1342_/B1 VDD VSS sg13g2_buf_1
XFILLER_62_393 VDD VSS sg13g2_decap_8
XFILLER_22_224 VDD VSS sg13g2_decap_8
XFILLER_50_511 VDD VSS sg13g2_decap_8
Xfanout39 fanout40/X _1338_/A2 VDD VSS sg13g2_buf_1
XFILLER_50_588 VDD VSS sg13g2_decap_4
XFILLER_109_819 VDD VSS sg13g2_decap_8
XFILLER_31_791 VDD VSS sg13g2_decap_8
XFILLER_13_49 VDD VSS sg13g2_decap_8
Xhold420 _2216_/Q VDD VSS _1383_/A sg13g2_dlygate4sd3_1
X_1829_ _1854_/A _1829_/A _2209_/Q VDD VSS sg13g2_nand2_1
Xhold453 _2303_/Q VDD VSS hold453/X sg13g2_dlygate4sd3_1
Xhold431 _2228_/Q VDD VSS _1414_/A sg13g2_dlygate4sd3_1
Xhold442 _1251_/Y VDD VSS _2357_/D sg13g2_dlygate4sd3_1
XFILLER_78_909 VDD VSS sg13g2_decap_8
XFILLER_104_524 VDD VSS sg13g2_decap_8
Xhold486 _2218_/Q VDD VSS _1389_/A sg13g2_dlygate4sd3_1
Xhold475 _2276_/Q VDD VSS hold475/X sg13g2_dlygate4sd3_1
Xhold464 _1568_/Y VDD VSS _1569_/B sg13g2_dlygate4sd3_1
XFILLER_89_279 VDD VSS sg13g2_decap_8
XFILLER_77_419 VDD VSS sg13g2_decap_8
Xhold497 _2274_/Q VDD VSS _1589_/A sg13g2_dlygate4sd3_1
XFILLER_38_35 VDD VSS sg13g2_decap_8
XFILLER_85_430 VDD VSS sg13g2_fill_2
XFILLER_58_644 VDD VSS sg13g2_decap_8
XFILLER_46_817 VDD VSS sg13g2_decap_8
XFILLER_57_143 VDD VSS sg13g2_decap_8
XFILLER_85_496 VDD VSS sg13g2_decap_8
XFILLER_54_850 VDD VSS sg13g2_decap_8
XFILLER_54_23 VDD VSS sg13g2_fill_1
XFILLER_38_390 VDD VSS sg13g2_decap_8
XFILLER_72_168 VDD VSS sg13g2_decap_8
XFILLER_26_574 VDD VSS sg13g2_decap_8
XFILLER_14_714 VDD VSS sg13g2_decap_8
XFILLER_81_680 VDD VSS sg13g2_decap_8
XFILLER_53_382 VDD VSS sg13g2_decap_8
XFILLER_13_224 VDD VSS sg13g2_decap_8
XFILLER_54_78 VDD VSS sg13g2_decap_8
XFILLER_110_84 VDD VSS sg13g2_decap_8
XFILLER_9_217 VDD VSS sg13g2_decap_8
XFILLER_16_1022 VDD VSS sg13g2_decap_8
XFILLER_70_77 VDD VSS sg13g2_decap_8
XFILLER_22_791 VDD VSS sg13g2_decap_8
XFILLER_10_931 VDD VSS sg13g2_decap_8
XFILLER_103_1036 VDD VSS sg13g2_decap_8
XFILLER_6_924 VDD VSS sg13g2_decap_8
XFILLER_5_434 VDD VSS sg13g2_decap_8
XFILLER_108_885 VDD VSS sg13g2_decap_8
XFILLER_79_42 VDD VSS sg13g2_decap_8
XFILLER_107_395 VDD VSS sg13g2_decap_8
XFILLER_96_728 VDD VSS sg13g2_decap_8
XFILLER_1_651 VDD VSS sg13g2_decap_8
XFILLER_49_622 VDD VSS sg13g2_decap_8
XFILLER_0_161 VDD VSS sg13g2_decap_8
XFILLER_88_290 VDD VSS sg13g2_decap_8
XFILLER_76_441 VDD VSS sg13g2_decap_8
XFILLER_95_63 VDD VSS sg13g2_decap_8
XFILLER_23_1015 VDD VSS sg13g2_decap_8
XFILLER_49_655 VDD VSS sg13g2_decap_8
XFILLER_48_132 VDD VSS sg13g2_decap_8
XFILLER_77_986 VDD VSS sg13g2_decap_8
XFILLER_48_154 VDD VSS sg13g2_fill_2
XFILLER_92_967 VDD VSS sg13g2_decap_8
XFILLER_91_433 VDD VSS sg13g2_decap_8
XFILLER_64_669 VDD VSS sg13g2_decap_8
XFILLER_51_319 VDD VSS sg13g2_decap_8
XFILLER_17_574 VDD VSS sg13g2_decap_8
XFILLER_60_820 VDD VSS sg13g2_decap_8
XFILLER_32_511 VDD VSS sg13g2_decap_8
XFILLER_44_371 VDD VSS sg13g2_decap_8
XFILLER_71_190 VDD VSS sg13g2_fill_2
XFILLER_60_886 VDD VSS sg13g2_decap_8
XFILLER_32_588 VDD VSS sg13g2_decap_8
XFILLER_20_728 VDD VSS sg13g2_decap_8
XFILLER_30_1008 VDD VSS sg13g2_decap_8
XFILLER_13_791 VDD VSS sg13g2_decap_8
XFILLER_9_784 VDD VSS sg13g2_decap_8
XFILLER_8_294 VDD VSS sg13g2_decap_8
X_1614_ _1613_/Y VDD _1614_/Y VSS _1638_/S hold547/X sg13g2_o21ai_1
XFILLER_99_555 VDD VSS sg13g2_decap_8
X_1545_ _1544_/Y VDD _1545_/Y VSS _1580_/A1 _2205_/Q sg13g2_o21ai_1
XFILLER_87_717 VDD VSS sg13g2_decap_8
XFILLER_101_527 VDD VSS sg13g2_decap_8
XFILLER_86_216 VDD VSS sg13g2_decap_8
X_1476_ _1602_/B VDD _1476_/Y VSS _1382_/A _1479_/A2 sg13g2_o21ai_1
XFILLER_95_794 VDD VSS sg13g2_decap_8
XFILLER_39_154 VDD VSS sg13g2_decap_8
XFILLER_83_967 VDD VSS sg13g2_decap_8
X_2200__140 VDD VSS _2200_/RESET_B sg13g2_tiehi
XFILLER_82_422 VDD VSS sg13g2_decap_8
XFILLER_55_669 VDD VSS sg13g2_decap_8
XFILLER_54_113 VDD VSS sg13g2_decap_8
XFILLER_78_1060 VDD VSS sg13g2_fill_1
X_2028_ _2027_/X _2074_/A _2025_/Y _2324_/D VDD VSS sg13g2_a21o_1
XFILLER_39_1011 VDD VSS sg13g2_decap_8
XFILLER_36_861 VDD VSS sg13g2_decap_8
XFILLER_54_168 VDD VSS sg13g2_decap_8
XFILLER_42_308 VDD VSS sg13g2_decap_4
XFILLER_82_499 VDD VSS sg13g2_decap_8
XFILLER_23_511 VDD VSS sg13g2_decap_8
XFILLER_35_371 VDD VSS sg13g2_decap_8
XFILLER_51_897 VDD VSS sg13g2_decap_8
XFILLER_23_588 VDD VSS sg13g2_decap_8
XFILLER_11_728 VDD VSS sg13g2_decap_8
XFILLER_50_374 VDD VSS sg13g2_decap_8
XFILLER_10_238 VDD VSS sg13g2_decap_8
XFILLER_109_616 VDD VSS sg13g2_decap_8
XFILLER_40_14 VDD VSS sg13g2_decap_8
XFILLER_108_126 VDD VSS sg13g2_decap_8
XFILLER_3_938 VDD VSS sg13g2_decap_8
XFILLER_105_833 VDD VSS sg13g2_decap_8
XFILLER_104_321 VDD VSS sg13g2_decap_8
XFILLER_2_448 VDD VSS sg13g2_decap_8
Xhold294 _1227_/Y VDD VSS _1228_/B sg13g2_dlygate4sd3_1
XFILLER_46_1059 VDD VSS sg13g2_fill_2
XFILLER_49_56 VDD VSS sg13g2_decap_8
XFILLER_77_249 VDD VSS sg13g2_decap_8
XFILLER_59_964 VDD VSS sg13g2_decap_8
XFILLER_58_452 VDD VSS sg13g2_fill_1
XFILLER_100_560 VDD VSS sg13g2_decap_8
XFILLER_74_912 VDD VSS sg13g2_decap_8
XFILLER_73_400 VDD VSS sg13g2_decap_8
XFILLER_105_84 VDD VSS sg13g2_decap_8
XFILLER_46_614 VDD VSS sg13g2_decap_8
XFILLER_73_477 VDD VSS sg13g2_decap_8
XFILLER_27_861 VDD VSS sg13g2_decap_8
XFILLER_45_146 VDD VSS sg13g2_decap_4
XFILLER_33_308 VDD VSS sg13g2_decap_8
XFILLER_45_168 VDD VSS sg13g2_decap_8
XFILLER_14_511 VDD VSS sg13g2_decap_8
XFILLER_26_371 VDD VSS sg13g2_decap_8
XFILLER_81_21 VDD VSS sg13g2_decap_8
XFILLER_42_875 VDD VSS sg13g2_decap_8
XFILLER_14_588 VDD VSS sg13g2_decap_8
XFILLER_81_98 VDD VSS sg13g2_decap_8
XFILLER_14_70 VDD VSS sg13g2_decap_8
XFILLER_6_721 VDD VSS sg13g2_decap_8
XFILLER_5_231 VDD VSS sg13g2_decap_8
XFILLER_108_682 VDD VSS sg13g2_decap_8
XFILLER_6_798 VDD VSS sg13g2_decap_8
XFILLER_30_91 VDD VSS sg13g2_decap_8
XFILLER_46_7 VDD VSS sg13g2_decap_8
XFILLER_69_706 VDD VSS sg13g2_decap_8
X_1330_ _1330_/Y _1482_/B1 hold404/X _1482_/A2 _2328_/Q VDD VSS sg13g2_a22oi_1
XFILLER_111_847 VDD VSS sg13g2_decap_8
X_2182__176 VDD VSS _2182_/RESET_B sg13g2_tiehi
XFILLER_96_514 VDD VSS sg13g2_decap_8
X_1261_ _2150_/A VDD _1261_/Y VSS _1255_/B _1516_/A sg13g2_o21ai_1
XFILLER_110_368 VDD VSS sg13g2_decap_8
XFILLER_65_923 VDD VSS sg13g2_decap_8
X_1192_ VDD _1492_/A _1192_/A VSS sg13g2_inv_1
XFILLER_49_485 VDD VSS sg13g2_decap_4
XFILLER_92_742 VDD VSS sg13g2_decap_8
XFILLER_76_282 VDD VSS sg13g2_decap_8
XFILLER_37_658 VDD VSS sg13g2_decap_8
XFILLER_91_241 VDD VSS sg13g2_decap_8
XFILLER_52_617 VDD VSS sg13g2_decap_8
XFILLER_18_861 VDD VSS sg13g2_decap_8
XFILLER_24_308 VDD VSS sg13g2_decap_8
XFILLER_36_168 VDD VSS sg13g2_decap_8
XFILLER_80_959 VDD VSS sg13g2_decap_8
XFILLER_17_371 VDD VSS sg13g2_decap_8
XFILLER_51_105 VDD VSS sg13g2_decap_8
XFILLER_33_875 VDD VSS sg13g2_decap_8
XFILLER_20_525 VDD VSS sg13g2_decap_8
XFILLER_32_385 VDD VSS sg13g2_decap_8
XFILLER_72_0 VDD VSS sg13g2_decap_8
XFILLER_9_581 VDD VSS sg13g2_decap_8
XFILLER_69_1059 VDD VSS sg13g2_fill_2
XFILLER_106_608 VDD VSS sg13g2_decap_8
XFILLER_10_28 VDD VSS sg13g2_decap_8
X_2341__139 VDD VSS _2341_/RESET_B sg13g2_tiehi
XFILLER_102_825 VDD VSS sg13g2_decap_8
XFILLER_101_302 VDD VSS sg13g2_decap_8
XFILLER_87_525 VDD VSS sg13g2_fill_2
XFILLER_87_514 VDD VSS sg13g2_decap_8
X_1528_ _1556_/S0 _2235_/Q _2227_/Q _2219_/Q _2211_/Q _1589_/B _1529_/A VDD VSS sg13g2_mux4_1
XFILLER_87_569 VDD VSS sg13g2_decap_8
XFILLER_68_750 VDD VSS sg13g2_decap_8
X_1459_ _1459_/A _1463_/B _1459_/Y VDD VSS sg13g2_nor2_1
XFILLER_101_379 VDD VSS sg13g2_decap_8
XFILLER_56_934 VDD VSS sg13g2_decap_8
XFILLER_28_658 VDD VSS sg13g2_decap_8
XFILLER_55_466 VDD VSS sg13g2_decap_8
XFILLER_15_308 VDD VSS sg13g2_decap_8
XFILLER_35_14 VDD VSS sg13g2_decap_8
XFILLER_27_168 VDD VSS sg13g2_decap_8
XFILLER_82_285 VDD VSS sg13g2_decap_8
XFILLER_70_414 VDD VSS sg13g2_decap_8
XFILLER_43_639 VDD VSS sg13g2_decap_8
XFILLER_42_105 VDD VSS sg13g2_decap_8
XFILLER_51_661 VDD VSS sg13g2_decap_8
XFILLER_24_875 VDD VSS sg13g2_decap_8
XFILLER_11_525 VDD VSS sg13g2_decap_8
XFILLER_23_385 VDD VSS sg13g2_decap_8
XFILLER_109_413 VDD VSS sg13g2_decap_8
XFILLER_52_1052 VDD VSS sg13g2_decap_8
XFILLER_7_518 VDD VSS sg13g2_decap_8
XFILLER_13_1036 VDD VSS sg13g2_decap_8
XFILLER_105_630 VDD VSS sg13g2_decap_8
XFILLER_3_735 VDD VSS sg13g2_decap_8
XFILLER_104_140 VDD VSS sg13g2_decap_8
XFILLER_2_245 VDD VSS sg13g2_decap_8
XFILLER_78_536 VDD VSS sg13g2_decap_4
XFILLER_104_195 VDD VSS sg13g2_decap_8
XFILLER_76_21 VDD VSS sg13g2_decap_8
XFILLER_59_772 VDD VSS sg13g2_fill_1
XFILLER_47_901 VDD VSS sg13g2_decap_4
XFILLER_65_219 VDD VSS sg13g2_decap_8
XFILLER_46_400 VDD VSS sg13g2_decap_8
XFILLER_86_591 VDD VSS sg13g2_decap_8
XFILLER_76_98 VDD VSS sg13g2_decap_8
XFILLER_19_658 VDD VSS sg13g2_decap_8
XFILLER_20_1029 VDD VSS sg13g2_decap_8
XFILLER_74_786 VDD VSS sg13g2_decap_8
XFILLER_100_390 VDD VSS sg13g2_fill_1
XFILLER_47_978 VDD VSS sg13g2_decap_8
XFILLER_18_168 VDD VSS sg13g2_decap_8
XFILLER_73_263 VDD VSS sg13g2_decap_8
XFILLER_92_42 VDD VSS sg13g2_decap_8
XFILLER_61_425 VDD VSS sg13g2_decap_8
XFILLER_33_105 VDD VSS sg13g2_decap_8
XFILLER_42_672 VDD VSS sg13g2_decap_8
XFILLER_30_812 VDD VSS sg13g2_decap_8
XFILLER_15_875 VDD VSS sg13g2_decap_8
XFILLER_14_385 VDD VSS sg13g2_decap_8
XFILLER_25_91 VDD VSS sg13g2_decap_8
XFILLER_30_889 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_3_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_109_980 VDD VSS sg13g2_decap_8
XFILLER_6_595 VDD VSS sg13g2_decap_8
XFILLER_29_1043 VDD VSS sg13g2_decap_8
X_2362_ _2362_/RESET_B VSS VDD _2362_/D _2362_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_111_644 VDD VSS sg13g2_decap_8
XFILLER_97_867 VDD VSS sg13g2_decap_8
XFILLER_69_558 VDD VSS sg13g2_decap_8
XFILLER_96_322 VDD VSS sg13g2_decap_8
X_1313_ VDD _2186_/D _1313_/A VSS sg13g2_inv_1
XFILLER_57_709 VDD VSS sg13g2_decap_8
X_2293_ _2293_/RESET_B VSS VDD _2293_/D _2293_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_84_517 VDD VSS sg13g2_fill_1
XFILLER_110_154 VDD VSS sg13g2_decap_8
XFILLER_38_912 VDD VSS sg13g2_decap_8
X_1244_ _1247_/C _2296_/Q _2258_/Q VDD VSS sg13g2_xnor2_1
XFILLER_49_260 VDD VSS sg13g2_decap_8
XFILLER_96_399 VDD VSS sg13g2_decap_8
XFILLER_65_731 VDD VSS sg13g2_fill_1
XFILLER_2_84 VDD VSS sg13g2_decap_8
XFILLER_38_989 VDD VSS sg13g2_decap_8
XFILLER_53_904 VDD VSS sg13g2_decap_8
XFILLER_37_455 VDD VSS sg13g2_decap_8
XFILLER_92_572 VDD VSS sg13g2_decap_8
XFILLER_53_937 VDD VSS sg13g2_fill_2
XFILLER_52_403 VDD VSS sg13g2_decap_8
XFILLER_24_105 VDD VSS sg13g2_decap_8
XFILLER_80_767 VDD VSS sg13g2_decap_8
XFILLER_75_1052 VDD VSS sg13g2_decap_8
XFILLER_36_1036 VDD VSS sg13g2_decap_8
XFILLER_33_672 VDD VSS sg13g2_decap_8
XFILLER_21_812 VDD VSS sg13g2_decap_8
XFILLER_20_322 VDD VSS sg13g2_decap_8
XFILLER_32_182 VDD VSS sg13g2_decap_8
XFILLER_21_889 VDD VSS sg13g2_decap_8
XFILLER_20_399 VDD VSS sg13g2_decap_8
XFILLER_21_49 VDD VSS sg13g2_decap_8
XFILLER_106_449 VDD VSS sg13g2_decap_8
XFILLER_82_1012 VDD VSS sg13g2_decap_8
XFILLER_88_823 VDD VSS sg13g2_decap_8
XFILLER_87_344 VDD VSS sg13g2_fill_1
XFILLER_0_749 VDD VSS sg13g2_decap_8
XFILLER_102_688 VDD VSS sg13g2_fill_1
XFILLER_102_677 VDD VSS sg13g2_fill_2
XFILLER_102_666 VDD VSS sg13g2_decap_8
XFILLER_87_388 VDD VSS sg13g2_decap_8
XFILLER_75_528 VDD VSS sg13g2_decap_8
XFILLER_101_198 VDD VSS sg13g2_decap_8
XFILLER_29_945 VDD VSS sg13g2_decap_8
XFILLER_56_742 VDD VSS sg13g2_decap_8
XFILLER_83_550 VDD VSS sg13g2_decap_8
XFILLER_55_252 VDD VSS sg13g2_decap_8
XFILLER_46_35 VDD VSS sg13g2_decap_8
XFILLER_28_455 VDD VSS sg13g2_decap_8
XFILLER_71_734 VDD VSS sg13g2_decap_8
XFILLER_15_105 VDD VSS sg13g2_decap_8
XFILLER_70_222 VDD VSS sg13g2_decap_8
XFILLER_102_63 VDD VSS sg13g2_decap_8
XFILLER_31_609 VDD VSS sg13g2_decap_8
X_2276__199 VDD VSS _2276_/RESET_B sg13g2_tiehi
XFILLER_70_255 VDD VSS sg13g2_decap_8
XFILLER_70_266 VDD VSS sg13g2_decap_8
XFILLER_24_672 VDD VSS sg13g2_decap_8
XFILLER_12_812 VDD VSS sg13g2_decap_8
XFILLER_30_119 VDD VSS sg13g2_decap_8
XFILLER_43_469 VDD VSS sg13g2_fill_2
XFILLER_70_299 VDD VSS sg13g2_decap_8
XFILLER_11_322 VDD VSS sg13g2_decap_8
XFILLER_8_805 VDD VSS sg13g2_decap_8
XFILLER_62_56 VDD VSS sg13g2_decap_8
XFILLER_23_182 VDD VSS sg13g2_decap_8
XFILLER_7_315 VDD VSS sg13g2_decap_8
XFILLER_12_889 VDD VSS sg13g2_decap_8
XFILLER_109_210 VDD VSS sg13g2_fill_2
XFILLER_11_399 VDD VSS sg13g2_decap_8
XFILLER_109_254 VDD VSS sg13g2_decap_8
XFILLER_3_532 VDD VSS sg13g2_decap_8
XFILLER_2_0 VDD VSS sg13g2_decap_8
XFILLER_106_972 VDD VSS sg13g2_decap_8
XFILLER_97_119 VDD VSS sg13g2_decap_8
XFILLER_87_42 VDD VSS sg13g2_decap_8
XFILLER_79_856 VDD VSS sg13g2_decap_4
XFILLER_93_303 VDD VSS sg13g2_decap_8
XFILLER_4_1001 VDD VSS sg13g2_decap_8
XFILLER_94_859 VDD VSS sg13g2_fill_2
XFILLER_93_369 VDD VSS sg13g2_decap_8
XFILLER_47_764 VDD VSS sg13g2_decap_8
XFILLER_19_455 VDD VSS sg13g2_decap_8
XFILLER_62_712 VDD VSS sg13g2_decap_8
XFILLER_46_263 VDD VSS sg13g2_decap_8
XFILLER_46_252 VDD VSS sg13g2_fill_2
XFILLER_35_959 VDD VSS sg13g2_decap_8
XFILLER_50_918 VDD VSS sg13g2_decap_8
XFILLER_62_789 VDD VSS sg13g2_fill_1
XFILLER_22_609 VDD VSS sg13g2_decap_8
XFILLER_61_266 VDD VSS sg13g2_decap_8
XFILLER_15_672 VDD VSS sg13g2_decap_8
XFILLER_34_469 VDD VSS sg13g2_decap_8
X_1931_ _1933_/B _1931_/A _1931_/B VDD VSS sg13g2_xnor2_1
XFILLER_14_182 VDD VSS sg13g2_decap_8
XFILLER_21_119 VDD VSS sg13g2_decap_8
X_1862_ _1862_/A _1852_/B _1863_/B VDD VSS sg13g2_nor2b_1
XFILLER_30_686 VDD VSS sg13g2_decap_8
X_1793_ _1795_/A _2216_/Q _2224_/Q VDD VSS sg13g2_nand2b_1
XFILLER_66_1007 VDD VSS sg13g2_decap_8
XFILLER_7_882 VDD VSS sg13g2_decap_8
XFILLER_6_392 VDD VSS sg13g2_decap_8
XFILLER_103_419 VDD VSS sg13g2_fill_2
XFILLER_88_119 VDD VSS sg13g2_decap_8
XFILLER_112_931 VDD VSS sg13g2_decap_8
XFILLER_35_0 VDD VSS sg13g2_decap_8
XFILLER_97_675 VDD VSS sg13g2_decap_8
X_2345_ _2345_/RESET_B VSS VDD _2345_/D _2345_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_111_441 VDD VSS sg13g2_decap_8
XFILLER_69_355 VDD VSS sg13g2_decap_8
XFILLER_69_366 VDD VSS sg13g2_fill_2
XFILLER_96_196 VDD VSS sg13g2_decap_8
X_2276_ _2276_/RESET_B VSS VDD _2276_/D _2276_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_57_528 VDD VSS sg13g2_decap_8
XFILLER_84_369 VDD VSS sg13g2_decap_8
XFILLER_65_550 VDD VSS sg13g2_decap_8
X_1227_ VSS VDD _1204_/Y _2365_/Q _1227_/Y _1500_/D sg13g2_a21oi_1
XFILLER_38_786 VDD VSS sg13g2_decap_8
XFILLER_37_252 VDD VSS sg13g2_decap_8
XFILLER_26_959 VDD VSS sg13g2_decap_8
XFILLER_16_49 VDD VSS sg13g2_decap_8
XFILLER_52_222 VDD VSS sg13g2_decap_4
XFILLER_13_609 VDD VSS sg13g2_decap_8
XFILLER_25_469 VDD VSS sg13g2_decap_8
XFILLER_12_119 VDD VSS sg13g2_decap_8
XFILLER_21_686 VDD VSS sg13g2_decap_8
XFILLER_20_196 VDD VSS sg13g2_decap_8
XFILLER_5_819 VDD VSS sg13g2_decap_8
XFILLER_106_224 VDD VSS sg13g2_decap_8
XFILLER_4_329 VDD VSS sg13g2_decap_8
XFILLER_107_758 VDD VSS sg13g2_decap_8
XFILLER_79_119 VDD VSS sg13g2_decap_8
XFILLER_103_931 VDD VSS sg13g2_decap_8
XFILLER_88_642 VDD VSS sg13g2_decap_8
XFILLER_0_546 VDD VSS sg13g2_decap_8
XFILLER_88_686 VDD VSS sg13g2_decap_8
XFILLER_76_804 VDD VSS sg13g2_fill_1
XFILLER_102_463 VDD VSS sg13g2_decap_8
XFILLER_87_130 VDD VSS sg13g2_decap_8
XFILLER_48_517 VDD VSS sg13g2_decap_4
XFILLER_76_837 VDD VSS sg13g2_decap_8
XFILLER_57_45 VDD VSS sg13g2_fill_1
XFILLER_57_67 VDD VSS sg13g2_decap_8
XFILLER_29_742 VDD VSS sg13g2_decap_8
XFILLER_84_892 VDD VSS sg13g2_decap_8
XFILLER_28_252 VDD VSS sg13g2_decap_8
XFILLER_44_767 VDD VSS sg13g2_decap_8
XFILLER_17_959 VDD VSS sg13g2_decap_8
XFILLER_71_564 VDD VSS sg13g2_decap_8
XFILLER_73_77 VDD VSS sg13g2_decap_8
XFILLER_16_469 VDD VSS sg13g2_decap_8
XFILLER_31_406 VDD VSS sg13g2_decap_8
XFILLER_43_244 VDD VSS sg13g2_decap_8
XFILLER_43_299 VDD VSS sg13g2_decap_8
XFILLER_8_602 VDD VSS sg13g2_decap_8
XFILLER_106_1056 VDD VSS sg13g2_decap_4
XFILLER_40_984 VDD VSS sg13g2_decap_8
XFILLER_7_112 VDD VSS sg13g2_decap_8
XFILLER_12_686 VDD VSS sg13g2_decap_8
XFILLER_89_1029 VDD VSS sg13g2_decap_8
XFILLER_11_196 VDD VSS sg13g2_decap_8
XFILLER_8_679 VDD VSS sg13g2_decap_8
XFILLER_22_70 VDD VSS sg13g2_decap_8
X_2326__207 VDD VSS _2326_/RESET_B sg13g2_tiehi
XFILLER_7_189 VDD VSS sg13g2_decap_8
XFILLER_98_439 VDD VSS sg13g2_decap_8
XFILLER_98_63 VDD VSS sg13g2_decap_8
XFILLER_4_896 VDD VSS sg13g2_decap_8
XFILLER_79_631 VDD VSS sg13g2_decap_8
XFILLER_112_238 VDD VSS sg13g2_decap_8
XFILLER_94_601 VDD VSS sg13g2_decap_8
XFILLER_79_664 VDD VSS sg13g2_decap_8
XFILLER_26_1057 VDD VSS sg13g2_decap_4
XFILLER_39_506 VDD VSS sg13g2_decap_8
X_2130_ _1688_/B VDD _2131_/B VSS _2142_/A1 hold526/X sg13g2_o21ai_1
X_2307__83 VDD VSS _2307__83/L_HI sg13g2_tiehi
XFILLER_67_848 VDD VSS sg13g2_decap_4
XFILLER_66_336 VDD VSS sg13g2_decap_4
X_2061_ _2047_/X _2049_/X _2061_/S _2062_/B VDD VSS sg13g2_mux2_1
XFILLER_93_133 VDD VSS sg13g2_decap_8
XFILLER_54_509 VDD VSS sg13g2_decap_8
XFILLER_47_583 VDD VSS sg13g2_decap_4
XFILLER_19_252 VDD VSS sg13g2_decap_8
XFILLER_35_756 VDD VSS sg13g2_decap_8
XFILLER_22_406 VDD VSS sg13g2_decap_8
XFILLER_34_266 VDD VSS sg13g2_decap_8
XFILLER_72_1011 VDD VSS sg13g2_decap_8
XFILLER_90_895 VDD VSS sg13g2_decap_8
X_1914_ _1919_/A _1914_/A _1914_/B VDD VSS sg13g2_xnor2_1
XFILLER_31_973 VDD VSS sg13g2_decap_8
XFILLER_30_483 VDD VSS sg13g2_decap_8
X_1845_ VDD VSS _1843_/X _1844_/X _1860_/A _1212_/Y _1856_/A _2206_/Q sg13g2_a221oi_1
X_1776_ _1809_/A _1776_/A _2226_/Q VDD VSS sg13g2_nand2_1
XFILLER_104_717 VDD VSS sg13g2_fill_1
XFILLER_103_249 VDD VSS sg13g2_decap_8
XFILLER_69_141 VDD VSS sg13g2_decap_8
XFILLER_100_945 VDD VSS sg13g2_decap_8
XFILLER_69_163 VDD VSS sg13g2_decap_8
X_2328_ _2328_/RESET_B VSS VDD _2328_/D _2328_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_57_369 VDD VSS sg13g2_decap_8
XFILLER_57_347 VDD VSS sg13g2_fill_2
XFILLER_85_689 VDD VSS sg13g2_decap_8
XFILLER_84_177 VDD VSS sg13g2_decap_8
XFILLER_38_583 VDD VSS sg13g2_decap_8
X_2259_ _2259_/RESET_B VSS VDD _2259_/D _2259_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_26_756 VDD VSS sg13g2_decap_8
XFILLER_13_406 VDD VSS sg13g2_decap_8
XFILLER_43_14 VDD VSS sg13g2_decap_8
XFILLER_25_266 VDD VSS sg13g2_decap_8
XFILLER_80_383 VDD VSS sg13g2_decap_8
XFILLER_41_748 VDD VSS sg13g2_decap_8
XFILLER_40_203 VDD VSS sg13g2_decap_8
XFILLER_22_973 VDD VSS sg13g2_decap_8
X_2210__120 VDD VSS _2210_/RESET_B sg13g2_tiehi
XFILLER_21_483 VDD VSS sg13g2_decap_8
XFILLER_107_500 VDD VSS sg13g2_decap_8
XFILLER_5_616 VDD VSS sg13g2_decap_8
XFILLER_107_555 VDD VSS sg13g2_decap_8
XFILLER_49_1002 VDD VSS sg13g2_decap_4
XFILLER_4_126 VDD VSS sg13g2_decap_8
XFILLER_49_1035 VDD VSS sg13g2_decap_8
XFILLER_108_84 VDD VSS sg13g2_decap_8
XFILLER_1_833 VDD VSS sg13g2_decap_8
XFILLER_88_450 VDD VSS sg13g2_decap_8
XFILLER_49_804 VDD VSS sg13g2_decap_8
XFILLER_0_343 VDD VSS sg13g2_decap_8
XFILLER_76_678 VDD VSS sg13g2_decap_8
XFILLER_84_21 VDD VSS sg13g2_decap_8
XFILLER_75_133 VDD VSS sg13g2_decap_8
XFILLER_48_336 VDD VSS sg13g2_decap_8
XFILLER_91_637 VDD VSS sg13g2_decap_8
XFILLER_1_1015 VDD VSS sg13g2_decap_8
XFILLER_95_1022 VDD VSS sg13g2_decap_8
XFILLER_75_199 VDD VSS sg13g2_fill_1
XFILLER_84_98 VDD VSS sg13g2_decap_8
XFILLER_56_391 VDD VSS sg13g2_decap_8
XFILLER_17_756 VDD VSS sg13g2_decap_8
XFILLER_44_564 VDD VSS sg13g2_decap_8
XFILLER_16_266 VDD VSS sg13g2_decap_8
XFILLER_17_70 VDD VSS sg13g2_decap_8
XFILLER_31_203 VDD VSS sg13g2_decap_8
XFILLER_40_781 VDD VSS sg13g2_decap_8
XFILLER_13_973 VDD VSS sg13g2_decap_8
XFILLER_76_7 VDD VSS sg13g2_decap_8
XFILLER_12_483 VDD VSS sg13g2_decap_8
XFILLER_9_966 VDD VSS sg13g2_decap_8
XFILLER_33_91 VDD VSS sg13g2_decap_8
XFILLER_32_1050 VDD VSS sg13g2_decap_8
XFILLER_8_476 VDD VSS sg13g2_decap_8
X_1630_ _1630_/Y _1634_/A _1630_/B VDD VSS sg13g2_nand2_1
XFILLER_99_715 VDD VSS sg13g2_decap_8
X_1561_ _1561_/Y _1527_/Y _1560_/Y hold461/X _1190_/Y VDD VSS sg13g2_a22oi_1
XFILLER_98_225 VDD VSS sg13g2_decap_8
X_1492_ _1492_/A _1492_/B _1495_/C _1493_/B VDD VSS sg13g2_nor3_1
XFILLER_4_693 VDD VSS sg13g2_decap_8
XFILLER_95_910 VDD VSS sg13g2_decap_8
XFILLER_79_461 VDD VSS sg13g2_decap_8
X_2113_ VSS VDD _2124_/B _2109_/X _2115_/A _2112_/Y sg13g2_a21oi_1
XFILLER_67_656 VDD VSS sg13g2_decap_8
XFILLER_55_818 VDD VSS sg13g2_decap_8
X_2296__125 VDD VSS _2296_/RESET_B sg13g2_tiehi
XFILLER_66_133 VDD VSS sg13g2_fill_2
XFILLER_95_987 VDD VSS sg13g2_decap_8
XFILLER_82_604 VDD VSS sg13g2_decap_8
XFILLER_94_475 VDD VSS sg13g2_decap_8
XFILLER_48_870 VDD VSS sg13g2_decap_8
XFILLER_54_306 VDD VSS sg13g2_decap_8
X_2337__155 VDD VSS _2337_/RESET_B sg13g2_tiehi
X_2044_ _2045_/A _2082_/B _2148_/B _2149_/A _1826_/B VDD VSS sg13g2_a22oi_1
XFILLER_66_188 VDD VSS sg13g2_decap_8
XFILLER_35_553 VDD VSS sg13g2_decap_8
X_2192__156 VDD VSS _2192_/RESET_B sg13g2_tiehi
Xfanout29 _1391_/Y _1392_/B VDD VSS sg13g2_buf_1
XFILLER_63_895 VDD VSS sg13g2_decap_8
Xfanout18 fanout22/X _1344_/B1 VDD VSS sg13g2_buf_1
XFILLER_22_203 VDD VSS sg13g2_decap_8
XFILLER_50_567 VDD VSS sg13g2_decap_8
XFILLER_31_770 VDD VSS sg13g2_decap_8
XFILLER_13_28 VDD VSS sg13g2_decap_8
XFILLER_30_280 VDD VSS sg13g2_decap_8
XFILLER_108_319 VDD VSS sg13g2_decap_8
X_1828_ _1876_/A _1874_/A _1874_/B VDD VSS sg13g2_nand2_1
Xhold410 _1517_/Y VDD VSS _2272_/D sg13g2_dlygate4sd3_1
Xhold454 _1660_/Y VDD VSS _1661_/B sg13g2_dlygate4sd3_1
X_1759_ _1760_/A _1760_/B _1927_/A VDD VSS sg13g2_and2_1
Xhold432 _2215_/Q VDD VSS _1380_/A sg13g2_dlygate4sd3_1
Xhold443 _2213_/Q VDD VSS _1374_/A sg13g2_dlygate4sd3_1
Xhold421 _2208_/Q VDD VSS hold421/X sg13g2_dlygate4sd3_1
Xhold465 _2214_/Q VDD VSS _1377_/A sg13g2_dlygate4sd3_1
XFILLER_89_225 VDD VSS sg13g2_fill_1
XFILLER_89_214 VDD VSS sg13g2_decap_8
Xhold487 _1390_/Y VDD VSS _2218_/D sg13g2_dlygate4sd3_1
Xhold476 _1540_/Y VDD VSS _1541_/B sg13g2_dlygate4sd3_1
XFILLER_89_258 VDD VSS sg13g2_decap_8
Xhold498 _1587_/Y VDD VSS _2286_/D sg13g2_dlygate4sd3_1
XFILLER_98_792 VDD VSS sg13g2_fill_2
XFILLER_58_623 VDD VSS sg13g2_decap_8
XFILLER_38_14 VDD VSS sg13g2_decap_8
XFILLER_86_965 VDD VSS sg13g2_decap_8
XFILLER_100_731 VDD VSS sg13g2_decap_8
XFILLER_57_122 VDD VSS sg13g2_decap_8
XFILLER_100_786 VDD VSS sg13g2_decap_8
XFILLER_73_604 VDD VSS sg13g2_fill_2
XFILLER_85_475 VDD VSS sg13g2_decap_8
XFILLER_39_892 VDD VSS sg13g2_decap_8
XFILLER_72_147 VDD VSS sg13g2_decap_8
XFILLER_26_553 VDD VSS sg13g2_decap_8
XFILLER_54_57 VDD VSS sg13g2_fill_2
XFILLER_54_35 VDD VSS sg13g2_decap_8
XFILLER_13_203 VDD VSS sg13g2_decap_8
XFILLER_41_523 VDD VSS sg13g2_fill_2
XFILLER_41_534 VDD VSS sg13g2_decap_4
XFILLER_16_1001 VDD VSS sg13g2_decap_8
XFILLER_110_63 VDD VSS sg13g2_decap_8
XFILLER_22_770 VDD VSS sg13g2_decap_8
XFILLER_10_910 VDD VSS sg13g2_decap_8
XFILLER_103_1015 VDD VSS sg13g2_decap_8
XFILLER_70_56 VDD VSS sg13g2_decap_8
XFILLER_6_903 VDD VSS sg13g2_decap_8
XFILLER_21_280 VDD VSS sg13g2_decap_8
XFILLER_5_413 VDD VSS sg13g2_decap_8
XFILLER_10_987 VDD VSS sg13g2_decap_8
XFILLER_108_864 VDD VSS sg13g2_decap_8
X_2222__96 VDD VSS _2222__96/L_HI sg13g2_tiehi
XFILLER_102_0 VDD VSS sg13g2_decap_8
XFILLER_79_21 VDD VSS sg13g2_decap_8
XFILLER_96_707 VDD VSS sg13g2_decap_8
XFILLER_79_98 VDD VSS sg13g2_decap_8
XFILLER_62_1010 VDD VSS sg13g2_fill_2
XFILLER_1_630 VDD VSS sg13g2_decap_8
XFILLER_0_140 VDD VSS sg13g2_decap_8
XFILLER_77_965 VDD VSS sg13g2_decap_8
XFILLER_95_42 VDD VSS sg13g2_decap_8
XFILLER_48_111 VDD VSS sg13g2_decap_8
XFILLER_110_1019 VDD VSS sg13g2_decap_8
XFILLER_92_946 VDD VSS sg13g2_decap_8
XFILLER_64_648 VDD VSS sg13g2_decap_8
XFILLER_28_91 VDD VSS sg13g2_decap_8
XFILLER_63_125 VDD VSS sg13g2_fill_2
XFILLER_17_553 VDD VSS sg13g2_decap_8
XFILLER_44_350 VDD VSS sg13g2_decap_8
XFILLER_91_489 VDD VSS sg13g2_decap_8
XFILLER_60_865 VDD VSS sg13g2_decap_8
XFILLER_32_567 VDD VSS sg13g2_decap_8
XFILLER_20_707 VDD VSS sg13g2_decap_8
XFILLER_13_770 VDD VSS sg13g2_decap_8
XFILLER_12_280 VDD VSS sg13g2_decap_8
XFILLER_9_763 VDD VSS sg13g2_decap_8
XFILLER_8_273 VDD VSS sg13g2_decap_8
X_1613_ _1613_/Y _1638_/S _1613_/B VDD VSS sg13g2_nand2_1
XFILLER_99_534 VDD VSS sg13g2_decap_8
X_1544_ VSS VDD _1580_/A1 _1213_/Y _1544_/Y _1523_/B sg13g2_a21oi_1
XFILLER_5_980 VDD VSS sg13g2_decap_8
XFILLER_101_506 VDD VSS sg13g2_decap_8
XFILLER_4_490 VDD VSS sg13g2_decap_8
XFILLER_5_84 VDD VSS sg13g2_decap_8
XIO_FILL_IO_EAST_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_1475_ VSS VDD _1197_/Y _1479_/A2 _2256_/D _1474_/Y sg13g2_a21oi_1
Xout_data_pads\[6\].out_data_pad _2372_/Q IOVDD IOVSS out_data_PADs[6] VDD VSS sg13g2_IOPadOut30mA
XFILLER_39_133 VDD VSS sg13g2_decap_8
XFILLER_83_924 VDD VSS sg13g2_fill_2
XFILLER_95_773 VDD VSS sg13g2_decap_8
XFILLER_83_913 VDD VSS sg13g2_decap_8
XFILLER_94_261 VDD VSS sg13g2_decap_8
XFILLER_82_401 VDD VSS sg13g2_decap_8
XFILLER_68_998 VDD VSS sg13g2_fill_1
XFILLER_67_464 VDD VSS sg13g2_decap_8
XFILLER_55_648 VDD VSS sg13g2_decap_8
XFILLER_36_840 VDD VSS sg13g2_decap_8
XFILLER_67_497 VDD VSS sg13g2_fill_2
X_2027_ _2036_/S _1949_/A _1878_/B _1889_/A _1826_/B _2054_/S _2027_/X VDD VSS sg13g2_mux4_1
XFILLER_82_478 VDD VSS sg13g2_decap_8
XFILLER_35_350 VDD VSS sg13g2_decap_8
XFILLER_63_670 VDD VSS sg13g2_decap_8
XFILLER_51_821 VDD VSS sg13g2_decap_8
XFILLER_62_180 VDD VSS sg13g2_fill_2
XFILLER_11_707 VDD VSS sg13g2_decap_8
XFILLER_24_49 VDD VSS sg13g2_decap_8
XFILLER_23_567 VDD VSS sg13g2_decap_8
XFILLER_10_217 VDD VSS sg13g2_decap_8
XFILLER_108_105 VDD VSS sg13g2_decap_8
XFILLER_105_812 VDD VSS sg13g2_decap_8
XFILLER_3_917 VDD VSS sg13g2_decap_8
XFILLER_85_1043 VDD VSS sg13g2_decap_8
XFILLER_104_300 VDD VSS sg13g2_decap_8
XFILLER_2_427 VDD VSS sg13g2_decap_8
XFILLER_6_7 VDD VSS sg13g2_decap_8
XFILLER_105_889 VDD VSS sg13g2_decap_8
XFILLER_78_718 VDD VSS sg13g2_decap_4
XFILLER_46_1038 VDD VSS sg13g2_decap_8
XFILLER_49_35 VDD VSS sg13g2_decap_8
Xhold295 _2268_/Q VDD VSS hold295/X sg13g2_dlygate4sd3_1
XFILLER_104_388 VDD VSS sg13g2_fill_2
XFILLER_104_377 VDD VSS sg13g2_decap_8
XFILLER_77_228 VDD VSS sg13g2_decap_8
XFILLER_49_79 VDD VSS sg13g2_decap_8
XFILLER_59_943 VDD VSS sg13g2_decap_8
XFILLER_105_63 VDD VSS sg13g2_decap_8
XFILLER_74_968 VDD VSS sg13g2_decap_8
XFILLER_86_795 VDD VSS sg13g2_decap_8
XFILLER_58_497 VDD VSS sg13g2_decap_8
XFILLER_45_125 VDD VSS sg13g2_decap_8
XFILLER_65_56 VDD VSS sg13g2_decap_8
XFILLER_73_456 VDD VSS sg13g2_decap_8
XFILLER_61_618 VDD VSS sg13g2_decap_8
XFILLER_27_840 VDD VSS sg13g2_decap_8
XFILLER_92_1025 VDD VSS sg13g2_fill_1
XFILLER_61_629 VDD VSS sg13g2_fill_1
XFILLER_54_670 VDD VSS sg13g2_fill_1
XFILLER_60_106 VDD VSS sg13g2_decap_8
XFILLER_26_350 VDD VSS sg13g2_decap_8
XFILLER_42_854 VDD VSS sg13g2_decap_8
XFILLER_81_77 VDD VSS sg13g2_decap_8
XFILLER_14_567 VDD VSS sg13g2_decap_8
XFILLER_6_700 VDD VSS sg13g2_decap_8
XFILLER_5_210 VDD VSS sg13g2_decap_8
XFILLER_10_784 VDD VSS sg13g2_decap_8
XFILLER_108_661 VDD VSS sg13g2_decap_8
XFILLER_6_777 VDD VSS sg13g2_decap_8
XFILLER_107_182 VDD VSS sg13g2_fill_1
XFILLER_5_287 VDD VSS sg13g2_decap_8
XFILLER_30_70 VDD VSS sg13g2_decap_8
XFILLER_107_193 VDD VSS sg13g2_decap_4
XFILLER_111_826 VDD VSS sg13g2_decap_8
XFILLER_2_994 VDD VSS sg13g2_decap_8
XFILLER_39_7 VDD VSS sg13g2_decap_8
XFILLER_110_347 VDD VSS sg13g2_decap_8
X_1260_ VSS VDD _1516_/A _1514_/A _1260_/A sg13g2_or2_1
XFILLER_68_239 VDD VSS sg13g2_decap_8
XFILLER_7_1043 VDD VSS sg13g2_decap_8
XFILLER_76_261 VDD VSS sg13g2_decap_8
XFILLER_65_902 VDD VSS sg13g2_decap_8
X_1191_ VDD _1366_/A _2267_/Q VSS sg13g2_inv_1
XFILLER_92_721 VDD VSS sg13g2_decap_8
XFILLER_77_795 VDD VSS sg13g2_decap_8
XFILLER_91_220 VDD VSS sg13g2_decap_8
XFILLER_37_637 VDD VSS sg13g2_decap_8
XFILLER_65_979 VDD VSS sg13g2_decap_8
XFILLER_18_840 VDD VSS sg13g2_decap_8
XFILLER_36_147 VDD VSS sg13g2_decap_8
XFILLER_92_798 VDD VSS sg13g2_decap_8
XFILLER_17_350 VDD VSS sg13g2_decap_8
XFILLER_33_854 VDD VSS sg13g2_decap_8
XFILLER_20_504 VDD VSS sg13g2_decap_8
XFILLER_32_364 VDD VSS sg13g2_decap_8
XFILLER_9_560 VDD VSS sg13g2_decap_8
XFILLER_65_0 VDD VSS sg13g2_decap_8
Xrst_n_pad IOVDD IOVSS fanout78/A rst_n_PAD VDD VSS sg13g2_IOPadIn
XFILLER_105_119 VDD VSS sg13g2_decap_8
XFILLER_99_353 VDD VSS sg13g2_decap_8
X_1527_ _1594_/A _1527_/B _1527_/Y VDD VSS sg13g2_nor2_1
XFILLER_87_548 VDD VSS sg13g2_decap_8
X_1458_ VSS VDD _1379_/Y _1463_/B _2248_/D _1457_/Y sg13g2_a21oi_1
XFILLER_101_358 VDD VSS sg13g2_decap_8
XFILLER_74_209 VDD VSS sg13g2_decap_8
XFILLER_56_913 VDD VSS sg13g2_fill_1
XFILLER_19_49 VDD VSS sg13g2_decap_8
X_1389_ _1389_/Y _1389_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_68_795 VDD VSS sg13g2_fill_1
XFILLER_28_637 VDD VSS sg13g2_decap_8
XFILLER_67_294 VDD VSS sg13g2_decap_8
XFILLER_55_445 VDD VSS sg13g2_decap_8
XFILLER_27_147 VDD VSS sg13g2_decap_8
XFILLER_71_949 VDD VSS sg13g2_decap_8
XFILLER_83_787 VDD VSS sg13g2_decap_8
XFILLER_82_264 VDD VSS sg13g2_decap_8
XFILLER_43_618 VDD VSS sg13g2_decap_8
XFILLER_51_640 VDD VSS sg13g2_decap_8
XFILLER_24_854 VDD VSS sg13g2_decap_8
XFILLER_11_504 VDD VSS sg13g2_decap_8
XFILLER_23_364 VDD VSS sg13g2_decap_8
XFILLER_51_14 VDD VSS sg13g2_decap_8
XFILLER_13_1015 VDD VSS sg13g2_decap_8
XFILLER_100_1018 VDD VSS sg13g2_decap_8
XFILLER_109_469 VDD VSS sg13g2_decap_8
XFILLER_3_714 VDD VSS sg13g2_decap_8
XFILLER_2_224 VDD VSS sg13g2_decap_8
XFILLER_105_686 VDD VSS sg13g2_decap_8
XFILLER_104_174 VDD VSS sg13g2_decap_8
XFILLER_78_515 VDD VSS sg13g2_decap_8
XFILLER_86_570 VDD VSS sg13g2_decap_8
XFILLER_76_77 VDD VSS sg13g2_decap_8
XFILLER_47_957 VDD VSS sg13g2_decap_8
XFILLER_19_637 VDD VSS sg13g2_decap_8
XFILLER_20_1008 VDD VSS sg13g2_decap_8
XFILLER_92_21 VDD VSS sg13g2_decap_8
XFILLER_18_147 VDD VSS sg13g2_decap_8
XFILLER_61_404 VDD VSS sg13g2_decap_8
XFILLER_46_489 VDD VSS sg13g2_decap_8
XFILLER_15_854 VDD VSS sg13g2_decap_8
XFILLER_109_1043 VDD VSS sg13g2_decap_8
XFILLER_92_98 VDD VSS sg13g2_decap_8
XFILLER_42_651 VDD VSS sg13g2_decap_8
XFILLER_14_364 VDD VSS sg13g2_decap_8
XFILLER_25_70 VDD VSS sg13g2_decap_8
XFILLER_30_868 VDD VSS sg13g2_decap_8
XFILLER_10_581 VDD VSS sg13g2_decap_8
XFILLER_41_91 VDD VSS sg13g2_decap_8
XFILLER_6_574 VDD VSS sg13g2_decap_8
XFILLER_29_1022 VDD VSS sg13g2_decap_8
XFILLER_96_301 VDD VSS sg13g2_decap_8
X_2361_ _2361_/RESET_B VSS VDD _2361_/D _2361_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_111_623 VDD VSS sg13g2_decap_8
XFILLER_97_846 VDD VSS sg13g2_decap_8
XFILLER_69_537 VDD VSS sg13g2_decap_8
X_1312_ _1312_/Y _1344_/B1 hold327/X _1344_/A2 _2350_/Q VDD VSS sg13g2_a22oi_1
XFILLER_2_791 VDD VSS sg13g2_decap_8
X_2292_ _2292_/RESET_B VSS VDD _2292_/D _2292_/Q clkload3/A sg13g2_dfrbpq_1
XFILLER_96_378 VDD VSS sg13g2_decap_8
XFILLER_110_133 VDD VSS sg13g2_decap_8
X_1243_ _1247_/B _2290_/Q _2252_/Q VDD VSS sg13g2_xnor2_1
XFILLER_65_710 VDD VSS sg13g2_decap_8
XFILLER_2_63 VDD VSS sg13g2_decap_8
XFILLER_37_434 VDD VSS sg13g2_decap_8
XFILLER_92_551 VDD VSS sg13g2_decap_8
XFILLER_92_540 VDD VSS sg13g2_decap_4
XFILLER_38_968 VDD VSS sg13g2_decap_8
XFILLER_65_787 VDD VSS sg13g2_fill_1
XFILLER_64_275 VDD VSS sg13g2_decap_8
XFILLER_80_746 VDD VSS sg13g2_decap_8
XFILLER_36_1015 VDD VSS sg13g2_decap_8
XFILLER_33_651 VDD VSS sg13g2_decap_8
XFILLER_61_993 VDD VSS sg13g2_fill_2
XFILLER_60_470 VDD VSS sg13g2_decap_8
XFILLER_20_301 VDD VSS sg13g2_decap_8
XFILLER_32_161 VDD VSS sg13g2_decap_8
XFILLER_21_868 VDD VSS sg13g2_decap_8
XFILLER_20_378 VDD VSS sg13g2_decap_8
XFILLER_21_28 VDD VSS sg13g2_decap_8
XFILLER_106_428 VDD VSS sg13g2_decap_8
XFILLER_88_802 VDD VSS sg13g2_decap_8
XFILLER_0_728 VDD VSS sg13g2_decap_8
XFILLER_102_623 VDD VSS sg13g2_decap_8
XFILLER_88_879 VDD VSS sg13g2_decap_8
XFILLER_101_133 VDD VSS sg13g2_decap_8
XFILLER_29_924 VDD VSS sg13g2_decap_8
XFILLER_56_721 VDD VSS sg13g2_decap_8
XFILLER_46_14 VDD VSS sg13g2_decap_8
XFILLER_55_231 VDD VSS sg13g2_decap_8
XFILLER_28_434 VDD VSS sg13g2_decap_8
XFILLER_71_713 VDD VSS sg13g2_decap_8
XFILLER_44_949 VDD VSS sg13g2_decap_8
XFILLER_56_798 VDD VSS sg13g2_decap_8
XFILLER_102_42 VDD VSS sg13g2_decap_8
XFILLER_43_448 VDD VSS sg13g2_decap_8
XFILLER_70_278 VDD VSS sg13g2_decap_8
XFILLER_24_651 VDD VSS sg13g2_decap_8
XFILLER_62_35 VDD VSS sg13g2_decap_8
XFILLER_11_301 VDD VSS sg13g2_decap_8
XFILLER_23_161 VDD VSS sg13g2_decap_8
XFILLER_12_868 VDD VSS sg13g2_decap_8
XFILLER_11_378 VDD VSS sg13g2_decap_8
XFILLER_109_288 VDD VSS sg13g2_fill_1
XFILLER_3_511 VDD VSS sg13g2_decap_8
XFILLER_106_951 VDD VSS sg13g2_decap_8
XFILLER_79_835 VDD VSS sg13g2_decap_8
XFILLER_87_21 VDD VSS sg13g2_decap_8
XFILLER_3_588 VDD VSS sg13g2_decap_8
XFILLER_105_483 VDD VSS sg13g2_decap_8
XFILLER_87_98 VDD VSS sg13g2_decap_8
X_2220__100 VDD VSS _2220_/RESET_B sg13g2_tiehi
XFILLER_78_389 VDD VSS sg13g2_decap_8
XFILLER_98_1053 VDD VSS sg13g2_decap_8
XFILLER_93_348 VDD VSS sg13g2_decap_8
XFILLER_47_743 VDD VSS sg13g2_decap_8
XFILLER_19_434 VDD VSS sg13g2_decap_8
XFILLER_4_1057 VDD VSS sg13g2_decap_4
XFILLER_46_220 VDD VSS sg13g2_decap_8
XFILLER_35_938 VDD VSS sg13g2_decap_8
XFILLER_62_702 VDD VSS sg13g2_fill_1
XFILLER_59_1059 VDD VSS sg13g2_fill_2
XFILLER_59_1048 VDD VSS sg13g2_decap_8
XFILLER_62_768 VDD VSS sg13g2_decap_8
XFILLER_61_234 VDD VSS sg13g2_decap_8
XFILLER_36_91 VDD VSS sg13g2_decap_8
XFILLER_34_448 VDD VSS sg13g2_decap_8
XFILLER_43_982 VDD VSS sg13g2_decap_8
XFILLER_15_651 VDD VSS sg13g2_decap_8
X_1930_ _1931_/B _1930_/A _1999_/A VDD VSS sg13g2_nand2_1
XFILLER_14_161 VDD VSS sg13g2_decap_8
X_1861_ _1892_/A _1952_/A _1952_/B VDD VSS sg13g2_nand2_1
XFILLER_30_665 VDD VSS sg13g2_decap_8
X_1792_ _2224_/Q _2216_/Q _1792_/Y VDD VSS sg13g2_nor2b_1
XFILLER_7_861 VDD VSS sg13g2_decap_8
XFILLER_6_371 VDD VSS sg13g2_decap_8
XFILLER_112_910 VDD VSS sg13g2_decap_8
XFILLER_97_621 VDD VSS sg13g2_fill_2
XFILLER_111_420 VDD VSS sg13g2_decap_8
XFILLER_69_334 VDD VSS sg13g2_decap_8
XFILLER_69_323 VDD VSS sg13g2_decap_8
X_2344_ _2344_/RESET_B VSS VDD _2344_/D _2344_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_112_987 VDD VSS sg13g2_decap_8
XFILLER_97_654 VDD VSS sg13g2_decap_8
XFILLER_85_805 VDD VSS sg13g2_fill_1
XFILLER_57_507 VDD VSS sg13g2_decap_8
XFILLER_28_0 VDD VSS sg13g2_decap_8
XFILLER_111_497 VDD VSS sg13g2_decap_8
XFILLER_96_175 VDD VSS sg13g2_decap_8
X_2275_ _2275_/RESET_B VSS VDD _2275_/D _2275_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_84_348 VDD VSS sg13g2_decap_8
XFILLER_38_765 VDD VSS sg13g2_decap_8
XFILLER_37_231 VDD VSS sg13g2_decap_8
X_1226_ _1226_/X _1236_/C _1226_/B _2361_/Q VDD VSS sg13g2_and3_1
XFILLER_26_938 VDD VSS sg13g2_decap_8
XFILLER_16_28 VDD VSS sg13g2_decap_8
XFILLER_25_448 VDD VSS sg13g2_decap_8
XFILLER_52_267 VDD VSS sg13g2_decap_8
XFILLER_21_665 VDD VSS sg13g2_decap_8
XFILLER_20_175 VDD VSS sg13g2_decap_8
XFILLER_32_49 VDD VSS sg13g2_decap_8
X_2347__113 VDD VSS _2347_/RESET_B sg13g2_tiehi
XFILLER_107_737 VDD VSS sg13g2_decap_8
XFILLER_106_203 VDD VSS sg13g2_decap_8
XFILLER_4_308 VDD VSS sg13g2_decap_8
XFILLER_10_1029 VDD VSS sg13g2_decap_8
XFILLER_106_7 VDD VSS sg13g2_decap_8
XFILLER_103_910 VDD VSS sg13g2_decap_8
XFILLER_88_621 VDD VSS sg13g2_decap_8
XFILLER_0_525 VDD VSS sg13g2_decap_8
XFILLER_103_987 VDD VSS sg13g2_decap_8
XFILLER_76_816 VDD VSS sg13g2_decap_8
XFILLER_102_442 VDD VSS sg13g2_decap_8
XFILLER_29_721 VDD VSS sg13g2_decap_8
XFILLER_91_808 VDD VSS sg13g2_decap_8
XFILLER_75_348 VDD VSS sg13g2_decap_8
XFILLER_28_231 VDD VSS sg13g2_decap_8
XFILLER_84_871 VDD VSS sg13g2_decap_8
XFILLER_29_798 VDD VSS sg13g2_decap_8
XFILLER_17_938 VDD VSS sg13g2_decap_8
XFILLER_71_543 VDD VSS sg13g2_decap_8
XFILLER_73_56 VDD VSS sg13g2_decap_8
XFILLER_56_595 VDD VSS sg13g2_decap_8
XFILLER_44_746 VDD VSS sg13g2_decap_8
XFILLER_16_448 VDD VSS sg13g2_decap_8
XFILLER_71_598 VDD VSS sg13g2_decap_8
XFILLER_19_1043 VDD VSS sg13g2_decap_8
XFILLER_106_1035 VDD VSS sg13g2_decap_8
XFILLER_40_963 VDD VSS sg13g2_decap_8
XFILLER_12_665 VDD VSS sg13g2_decap_8
XFILLER_11_175 VDD VSS sg13g2_decap_8
XFILLER_8_658 VDD VSS sg13g2_decap_8
XFILLER_7_168 VDD VSS sg13g2_decap_8
XFILLER_98_42 VDD VSS sg13g2_decap_8
XFILLER_79_610 VDD VSS sg13g2_decap_8
XFILLER_98_418 VDD VSS sg13g2_decap_8
XFILLER_4_875 VDD VSS sg13g2_decap_8
XFILLER_112_217 VDD VSS sg13g2_decap_8
XFILLER_3_385 VDD VSS sg13g2_decap_8
XFILLER_26_1036 VDD VSS sg13g2_decap_8
XFILLER_93_112 VDD VSS sg13g2_decap_8
XFILLER_67_827 VDD VSS sg13g2_decap_8
XFILLER_66_315 VDD VSS sg13g2_decap_8
XFILLER_21_7 VDD VSS sg13g2_decap_8
X_2060_ _2059_/Y VDD _2337_/D VSS _2025_/A _2055_/Y sg13g2_o21ai_1
XFILLER_19_231 VDD VSS sg13g2_decap_8
XFILLER_93_178 VDD VSS sg13g2_decap_8
XFILLER_47_595 VDD VSS sg13g2_fill_2
XFILLER_35_735 VDD VSS sg13g2_decap_8
XFILLER_62_554 VDD VSS sg13g2_decap_8
XFILLER_50_705 VDD VSS sg13g2_fill_1
XFILLER_34_245 VDD VSS sg13g2_decap_8
XFILLER_50_749 VDD VSS sg13g2_decap_8
X_1913_ _1930_/A VDD _1914_/B VSS _1816_/B _1901_/B sg13g2_o21ai_1
XFILLER_31_952 VDD VSS sg13g2_decap_8
XFILLER_33_1029 VDD VSS sg13g2_decap_8
XFILLER_30_462 VDD VSS sg13g2_decap_8
X_1844_ _1920_/A _1844_/B _1844_/X VDD VSS sg13g2_and2_1
XIO_FILL_IO_SOUTH_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_8_84 VDD VSS sg13g2_decap_8
X_1775_ _1874_/A _1775_/A _1775_/B VDD VSS sg13g2_xnor2_1
XFILLER_104_729 VDD VSS sg13g2_decap_8
XFILLER_69_120 VDD VSS sg13g2_decap_8
XFILLER_58_816 VDD VSS sg13g2_fill_1
XFILLER_112_784 VDD VSS sg13g2_decap_8
XFILLER_85_624 VDD VSS sg13g2_decap_8
X_2327_ _2327_/RESET_B VSS VDD _2327_/D _2327_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_84_112 VDD VSS sg13g2_decap_8
XFILLER_57_304 VDD VSS sg13g2_decap_8
XFILLER_85_668 VDD VSS sg13g2_decap_8
XFILLER_111_294 VDD VSS sg13g2_decap_8
XFILLER_57_337 VDD VSS sg13g2_fill_1
X_2258_ _2258_/RESET_B VSS VDD _2258_/D _2258_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_84_156 VDD VSS sg13g2_decap_8
XFILLER_38_562 VDD VSS sg13g2_decap_8
X_1209_ VDD _1829_/A _2250_/Q VSS sg13g2_inv_1
XFILLER_27_49 VDD VSS sg13g2_decap_8
X_2189_ _2189_/RESET_B VSS VDD _2189_/D _2189_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_66_893 VDD VSS sg13g2_decap_8
XFILLER_26_735 VDD VSS sg13g2_decap_8
XFILLER_65_392 VDD VSS sg13g2_decap_8
XFILLER_25_245 VDD VSS sg13g2_decap_8
XFILLER_80_362 VDD VSS sg13g2_decap_8
XFILLER_41_727 VDD VSS sg13g2_decap_8
XFILLER_22_952 VDD VSS sg13g2_decap_8
XFILLER_40_259 VDD VSS sg13g2_fill_1
XFILLER_21_462 VDD VSS sg13g2_decap_8
XFILLER_4_105 VDD VSS sg13g2_decap_8
XFILLER_107_534 VDD VSS sg13g2_decap_8
XFILLER_108_63 VDD VSS sg13g2_decap_8
XFILLER_1_812 VDD VSS sg13g2_decap_8
XFILLER_103_740 VDD VSS sg13g2_fill_2
XFILLER_0_322 VDD VSS sg13g2_decap_8
XFILLER_68_56 VDD VSS sg13g2_decap_4
XFILLER_89_996 VDD VSS sg13g2_decap_8
XFILLER_103_784 VDD VSS sg13g2_decap_8
XFILLER_75_112 VDD VSS sg13g2_decap_8
XFILLER_1_889 VDD VSS sg13g2_decap_8
XFILLER_68_89 VDD VSS sg13g2_decap_8
XFILLER_48_315 VDD VSS sg13g2_decap_8
XFILLER_76_657 VDD VSS sg13g2_decap_8
XFILLER_102_283 VDD VSS sg13g2_fill_1
XFILLER_102_294 VDD VSS sg13g2_decap_8
XFILLER_0_399 VDD VSS sg13g2_decap_8
XFILLER_48_359 VDD VSS sg13g2_fill_1
XFILLER_112_1050 VDD VSS sg13g2_decap_8
XFILLER_95_1001 VDD VSS sg13g2_decap_8
XFILLER_91_616 VDD VSS sg13g2_decap_8
XFILLER_75_178 VDD VSS sg13g2_decap_8
XFILLER_63_318 VDD VSS sg13g2_fill_2
XFILLER_84_690 VDD VSS sg13g2_decap_8
XFILLER_84_77 VDD VSS sg13g2_decap_8
XFILLER_29_595 VDD VSS sg13g2_decap_8
XFILLER_56_370 VDD VSS sg13g2_decap_8
XFILLER_17_735 VDD VSS sg13g2_decap_8
XFILLER_44_543 VDD VSS sg13g2_decap_8
XFILLER_16_245 VDD VSS sg13g2_decap_8
XFILLER_56_1029 VDD VSS sg13g2_decap_8
XFILLER_32_749 VDD VSS sg13g2_decap_8
XFILLER_13_952 VDD VSS sg13g2_decap_8
XFILLER_31_259 VDD VSS sg13g2_decap_8
XFILLER_40_760 VDD VSS sg13g2_decap_8
XFILLER_12_462 VDD VSS sg13g2_decap_8
XFILLER_9_945 VDD VSS sg13g2_decap_8
XFILLER_33_70 VDD VSS sg13g2_decap_8
XFILLER_8_455 VDD VSS sg13g2_decap_8
XFILLER_69_7 VDD VSS sg13g2_decap_8
X_1560_ _1559_/Y VDD _1560_/Y VSS _1592_/A _1557_/Y sg13g2_o21ai_1
XFILLER_98_204 VDD VSS sg13g2_decap_8
XFILLER_99_738 VDD VSS sg13g2_fill_1
X_1491_ _1495_/C _1497_/A _1491_/C _2265_/D VDD VSS sg13g2_nor3_1
XFILLER_4_672 VDD VSS sg13g2_decap_8
XFILLER_79_440 VDD VSS sg13g2_decap_8
XFILLER_3_182 VDD VSS sg13g2_decap_8
XFILLER_67_635 VDD VSS sg13g2_decap_8
XFILLER_95_966 VDD VSS sg13g2_decap_8
XFILLER_94_454 VDD VSS sg13g2_decap_8
X_2112_ _1259_/A VDD _2112_/Y VSS _2110_/Y _2111_/Y sg13g2_o21ai_1
XFILLER_66_112 VDD VSS sg13g2_decap_8
XFILLER_39_359 VDD VSS sg13g2_decap_8
XFILLER_66_167 VDD VSS sg13g2_decap_8
X_2043_ _2024_/X _2027_/X _2043_/S _2148_/B VDD VSS sg13g2_mux2_1
XFILLER_35_532 VDD VSS sg13g2_decap_8
XFILLER_47_392 VDD VSS sg13g2_decap_8
XFILLER_63_874 VDD VSS sg13g2_decap_8
XFILLER_62_351 VDD VSS sg13g2_decap_8
XFILLER_90_682 VDD VSS sg13g2_decap_8
Xfanout19 fanout22/X _1280_/B1 VDD VSS sg13g2_buf_1
XFILLER_23_749 VDD VSS sg13g2_decap_8
XFILLER_95_0 VDD VSS sg13g2_decap_8
XFILLER_50_546 VDD VSS sg13g2_decap_8
XFILLER_22_259 VDD VSS sg13g2_decap_8
X_2268__217 VDD VSS _2268_/RESET_B sg13g2_tiehi
X_1827_ VDD _1874_/B _1827_/A VSS sg13g2_inv_1
Xhold400 _1338_/Y VDD VSS _1339_/A sg13g2_dlygate4sd3_1
Xhold411 _2351_/Q VDD VSS _2099_/B sg13g2_dlygate4sd3_1
Xhold433 _2301_/Q VDD VSS _1697_/B sg13g2_dlygate4sd3_1
X_1758_ _1741_/Y VDD _1774_/B VSS _1772_/A _1772_/B sg13g2_o21ai_1
XIO_BOND_in_data_pads\[7\].in_data_pad in_data_PADs[7] bondpad_70x70
Xhold422 _2306_/Q VDD VSS hold422/X sg13g2_dlygate4sd3_1
X_2344__127 VDD VSS _2344_/RESET_B sg13g2_tiehi
Xhold444 _2249_/Q VDD VSS _1459_/A sg13g2_dlygate4sd3_1
XFILLER_2_609 VDD VSS sg13g2_decap_8
Xhold466 _2315_/Q VDD VSS hold466/X sg13g2_dlygate4sd3_1
Xhold477 _2238_/Q VDD VSS hold477/X sg13g2_dlygate4sd3_1
XFILLER_89_237 VDD VSS sg13g2_decap_8
X_1689_ _1687_/Y VDD _1689_/Y VSS _1724_/S hold490/X sg13g2_o21ai_1
Xhold455 _2206_/Q VDD VSS hold455/X sg13g2_dlygate4sd3_1
XFILLER_1_119 VDD VSS sg13g2_decap_8
Xhold488 _2204_/Q VDD VSS hold488/X sg13g2_dlygate4sd3_1
Xhold499 _2245_/Q VDD VSS _1451_/A sg13g2_dlygate4sd3_1
XFILLER_100_710 VDD VSS sg13g2_decap_8
XFILLER_98_771 VDD VSS sg13g2_decap_8
XFILLER_97_270 VDD VSS sg13g2_decap_8
XFILLER_86_944 VDD VSS sg13g2_decap_8
XFILLER_112_581 VDD VSS sg13g2_decap_8
XFILLER_100_754 VDD VSS sg13g2_fill_2
XFILLER_100_765 VDD VSS sg13g2_decap_8
XFILLER_73_616 VDD VSS sg13g2_decap_8
XFILLER_85_465 VDD VSS sg13g2_fill_2
XFILLER_85_454 VDD VSS sg13g2_decap_8
XFILLER_58_679 VDD VSS sg13g2_decap_8
XFILLER_39_871 VDD VSS sg13g2_decap_8
XFILLER_72_115 VDD VSS sg13g2_decap_4
XFILLER_54_14 VDD VSS sg13g2_decap_8
XFILLER_26_532 VDD VSS sg13g2_decap_8
XFILLER_45_329 VDD VSS sg13g2_decap_8
XFILLER_54_885 VDD VSS sg13g2_decap_8
XFILLER_41_502 VDD VSS sg13g2_decap_8
XFILLER_80_192 VDD VSS sg13g2_decap_8
XFILLER_110_42 VDD VSS sg13g2_decap_8
XFILLER_41_557 VDD VSS sg13g2_fill_2
XFILLER_14_749 VDD VSS sg13g2_decap_8
XFILLER_70_35 VDD VSS sg13g2_decap_8
XFILLER_13_259 VDD VSS sg13g2_decap_8
XFILLER_16_1057 VDD VSS sg13g2_decap_4
XFILLER_10_966 VDD VSS sg13g2_decap_8
XFILLER_108_843 VDD VSS sg13g2_decap_8
XFILLER_6_959 VDD VSS sg13g2_decap_8
XFILLER_107_353 VDD VSS sg13g2_decap_8
XFILLER_5_469 VDD VSS sg13g2_decap_8
XFILLER_79_77 VDD VSS sg13g2_decap_8
XFILLER_77_933 VDD VSS sg13g2_fill_2
XFILLER_110_529 VDD VSS sg13g2_decap_8
XFILLER_95_207 VDD VSS sg13g2_fill_1
XFILLER_95_21 VDD VSS sg13g2_decap_8
XFILLER_1_686 VDD VSS sg13g2_decap_8
XFILLER_103_581 VDD VSS sg13g2_decap_8
XFILLER_0_196 VDD VSS sg13g2_decap_8
XFILLER_76_476 VDD VSS sg13g2_decap_8
XFILLER_95_98 VDD VSS sg13g2_decap_8
XFILLER_64_627 VDD VSS sg13g2_decap_8
XFILLER_37_819 VDD VSS sg13g2_decap_8
XFILLER_48_156 VDD VSS sg13g2_fill_1
XFILLER_28_70 VDD VSS sg13g2_decap_8
XFILLER_63_104 VDD VSS sg13g2_decap_8
XFILLER_36_329 VDD VSS sg13g2_decap_8
XFILLER_48_189 VDD VSS sg13g2_decap_8
XFILLER_91_468 VDD VSS sg13g2_decap_8
XFILLER_17_532 VDD VSS sg13g2_decap_8
XFILLER_63_159 VDD VSS sg13g2_decap_8
XFILLER_29_392 VDD VSS sg13g2_decap_8
XFILLER_72_682 VDD VSS sg13g2_decap_8
XFILLER_71_192 VDD VSS sg13g2_fill_1
XFILLER_60_844 VDD VSS sg13g2_decap_8
XFILLER_32_546 VDD VSS sg13g2_decap_8
XFILLER_44_91 VDD VSS sg13g2_fill_2
XFILLER_9_742 VDD VSS sg13g2_decap_8
XFILLER_8_252 VDD VSS sg13g2_decap_8
X_1612_ _1613_/B _1612_/A _1617_/A VDD VSS sg13g2_xnor2_1
X_1543_ VDD _1543_/Y _1543_/A VSS sg13g2_inv_1
XFILLER_5_63 VDD VSS sg13g2_decap_8
X_1474_ _1602_/B VDD _1474_/Y VSS _1379_/A _1479_/A2 sg13g2_o21ai_1
XFILLER_68_911 VDD VSS sg13g2_decap_4
XFILLER_79_270 VDD VSS sg13g2_fill_1
XFILLER_68_966 VDD VSS sg13g2_fill_2
XFILLER_68_955 VDD VSS sg13g2_decap_8
XFILLER_67_443 VDD VSS sg13g2_decap_8
XFILLER_39_112 VDD VSS sg13g2_decap_8
XFILLER_94_240 VDD VSS sg13g2_decap_8
XFILLER_28_819 VDD VSS sg13g2_decap_8
XFILLER_10_0 VDD VSS sg13g2_decap_8
XFILLER_55_627 VDD VSS sg13g2_decap_8
XFILLER_27_329 VDD VSS sg13g2_decap_8
XFILLER_39_189 VDD VSS sg13g2_decap_8
X_2026_ _1878_/B _1826_/B _2054_/S _2026_/X VDD VSS sg13g2_mux2_1
XFILLER_70_619 VDD VSS sg13g2_decap_8
XFILLER_54_148 VDD VSS sg13g2_fill_2
XFILLER_39_1046 VDD VSS sg13g2_decap_8
XFILLER_51_800 VDD VSS sg13g2_decap_8
XFILLER_36_896 VDD VSS sg13g2_decap_8
XFILLER_90_490 VDD VSS sg13g2_decap_8
XFILLER_23_546 VDD VSS sg13g2_decap_8
XFILLER_62_192 VDD VSS sg13g2_decap_8
XFILLER_24_28 VDD VSS sg13g2_decap_8
XFILLER_50_332 VDD VSS sg13g2_decap_8
XFILLER_40_49 VDD VSS sg13g2_decap_8
XFILLER_2_406 VDD VSS sg13g2_decap_8
XFILLER_105_868 VDD VSS sg13g2_decap_8
XFILLER_104_356 VDD VSS sg13g2_decap_8
XFILLER_46_1017 VDD VSS sg13g2_decap_8
XFILLER_49_14 VDD VSS sg13g2_decap_8
Xhold296 _1499_/Y VDD VSS _2268_/D sg13g2_dlygate4sd3_1
X_2322__222 VDD VSS _2322_/RESET_B sg13g2_tiehi
XFILLER_59_922 VDD VSS sg13g2_decap_8
XFILLER_105_42 VDD VSS sg13g2_decap_8
X_2373__93 VDD VSS _2373__93/L_HI sg13g2_tiehi
XFILLER_58_443 VDD VSS sg13g2_decap_8
XFILLER_86_774 VDD VSS sg13g2_decap_8
XFILLER_59_999 VDD VSS sg13g2_decap_8
XFILLER_19_819 VDD VSS sg13g2_decap_8
XFILLER_74_947 VDD VSS sg13g2_decap_8
XFILLER_100_595 VDD VSS sg13g2_decap_8
XFILLER_85_273 VDD VSS sg13g2_decap_8
XFILLER_73_435 VDD VSS sg13g2_decap_8
XFILLER_22_1050 VDD VSS sg13g2_decap_8
XFILLER_46_638 VDD VSS sg13g2_decap_8
X_2279__187 VDD VSS _2279_/RESET_B sg13g2_tiehi
XFILLER_18_329 VDD VSS sg13g2_decap_8
XFILLER_65_35 VDD VSS sg13g2_decap_8
XFILLER_73_446 VDD VSS sg13g2_decap_4
XFILLER_82_991 VDD VSS sg13g2_decap_8
XFILLER_27_896 VDD VSS sg13g2_decap_8
XFILLER_42_833 VDD VSS sg13g2_decap_8
XFILLER_14_546 VDD VSS sg13g2_decap_8
XFILLER_81_56 VDD VSS sg13g2_decap_8
XFILLER_41_343 VDD VSS sg13g2_decap_8
XFILLER_10_763 VDD VSS sg13g2_decap_8
XFILLER_108_640 VDD VSS sg13g2_decap_8
XFILLER_6_756 VDD VSS sg13g2_decap_8
XFILLER_107_161 VDD VSS sg13g2_decap_8
XFILLER_5_266 VDD VSS sg13g2_decap_8
XFILLER_111_805 VDD VSS sg13g2_decap_8
XFILLER_68_218 VDD VSS sg13g2_decap_8
XFILLER_2_973 VDD VSS sg13g2_decap_8
XFILLER_110_326 VDD VSS sg13g2_decap_8
XFILLER_1_483 VDD VSS sg13g2_decap_8
XFILLER_7_1022 VDD VSS sg13g2_decap_8
XFILLER_77_774 VDD VSS sg13g2_decap_8
XFILLER_76_240 VDD VSS sg13g2_decap_8
XFILLER_37_616 VDD VSS sg13g2_decap_8
XFILLER_39_91 VDD VSS sg13g2_decap_8
X_1190_ VDD _1190_/Y _1589_/A VSS sg13g2_inv_1
XFILLER_49_454 VDD VSS sg13g2_decap_8
XFILLER_65_958 VDD VSS sg13g2_decap_8
XFILLER_64_402 VDD VSS sg13g2_decap_8
XFILLER_36_126 VDD VSS sg13g2_decap_8
XFILLER_92_777 VDD VSS sg13g2_decap_8
XFILLER_91_276 VDD VSS sg13g2_decap_4
XFILLER_64_479 VDD VSS sg13g2_decap_8
XFILLER_18_896 VDD VSS sg13g2_decap_8
XFILLER_72_490 VDD VSS sg13g2_decap_8
XFILLER_33_833 VDD VSS sg13g2_decap_8
XFILLER_60_652 VDD VSS sg13g2_fill_2
XFILLER_32_343 VDD VSS sg13g2_decap_8
XFILLER_69_1006 VDD VSS sg13g2_decap_8
XFILLER_58_0 VDD VSS sg13g2_decap_8
XFILLER_99_332 VDD VSS sg13g2_decap_8
X_1526_ _2284_/D _1524_/Y _2283_/D _2274_/D VDD VSS sg13g2_a21o_1
XFILLER_99_387 VDD VSS sg13g2_decap_8
XFILLER_101_337 VDD VSS sg13g2_decap_8
X_1457_ _1457_/A _1463_/B _1457_/Y VDD VSS sg13g2_nor2_1
XFILLER_59_229 VDD VSS sg13g2_decap_8
XFILLER_19_28 VDD VSS sg13g2_decap_8
X_1388_ _1388_/Y _1388_/A _1388_/B VDD VSS sg13g2_nand2_1
XFILLER_28_616 VDD VSS sg13g2_decap_8
XFILLER_67_251 VDD VSS sg13g2_decap_8
X_2370__85 VDD VSS _2370__85/L_HI sg13g2_tiehi
XFILLER_110_893 VDD VSS sg13g2_decap_8
XFILLER_95_582 VDD VSS sg13g2_decap_8
XFILLER_83_733 VDD VSS sg13g2_decap_8
XFILLER_68_785 VDD VSS sg13g2_decap_4
XFILLER_67_273 VDD VSS sg13g2_decap_8
XFILLER_55_424 VDD VSS sg13g2_decap_8
XFILLER_27_126 VDD VSS sg13g2_decap_8
XFILLER_83_766 VDD VSS sg13g2_decap_8
XFILLER_82_243 VDD VSS sg13g2_decap_8
XFILLER_71_928 VDD VSS sg13g2_decap_8
XFILLER_70_427 VDD VSS sg13g2_decap_4
XFILLER_35_49 VDD VSS sg13g2_decap_8
X_2009_ _1914_/A _1949_/A _2021_/S _2009_/X VDD VSS sg13g2_mux2_1
XFILLER_70_449 VDD VSS sg13g2_decap_8
XFILLER_36_693 VDD VSS sg13g2_decap_8
XFILLER_24_833 VDD VSS sg13g2_decap_8
XFILLER_50_151 VDD VSS sg13g2_decap_8
XFILLER_23_343 VDD VSS sg13g2_decap_8
XFILLER_51_696 VDD VSS sg13g2_decap_8
XFILLER_50_195 VDD VSS sg13g2_decap_8
XFILLER_109_448 VDD VSS sg13g2_decap_8
XFILLER_2_203 VDD VSS sg13g2_decap_8
X_2207__126 VDD VSS _2207_/RESET_B sg13g2_tiehi
XFILLER_105_665 VDD VSS sg13g2_decap_8
XFILLER_93_519 VDD VSS sg13g2_decap_8
XFILLER_76_56 VDD VSS sg13g2_decap_8
XFILLER_59_763 VDD VSS sg13g2_fill_1
XFILLER_100_370 VDD VSS sg13g2_fill_1
XFILLER_47_936 VDD VSS sg13g2_decap_8
XFILLER_59_796 VDD VSS sg13g2_decap_8
XFILLER_19_616 VDD VSS sg13g2_decap_8
XFILLER_74_755 VDD VSS sg13g2_decap_4
XFILLER_73_243 VDD VSS sg13g2_decap_8
XFILLER_62_906 VDD VSS sg13g2_fill_2
XFILLER_58_295 VDD VSS sg13g2_decap_8
XFILLER_18_126 VDD VSS sg13g2_decap_8
XFILLER_46_468 VDD VSS sg13g2_decap_8
XFILLER_62_939 VDD VSS sg13g2_decap_8
XFILLER_55_980 VDD VSS sg13g2_decap_8
XFILLER_92_77 VDD VSS sg13g2_decap_8
XFILLER_42_630 VDD VSS sg13g2_decap_8
XFILLER_27_693 VDD VSS sg13g2_decap_8
XFILLER_15_833 VDD VSS sg13g2_decap_8
XFILLER_109_1022 VDD VSS sg13g2_decap_8
XFILLER_70_983 VDD VSS sg13g2_decap_8
XFILLER_14_343 VDD VSS sg13g2_decap_8
XFILLER_41_140 VDD VSS sg13g2_decap_8
XFILLER_30_847 VDD VSS sg13g2_decap_8
XFILLER_41_195 VDD VSS sg13g2_decap_8
XFILLER_10_560 VDD VSS sg13g2_decap_8
XFILLER_6_553 VDD VSS sg13g2_decap_8
XFILLER_41_70 VDD VSS sg13g2_decap_8
XFILLER_51_7 VDD VSS sg13g2_decap_8
XFILLER_108_492 VDD VSS sg13g2_fill_1
XFILLER_29_1001 VDD VSS sg13g2_decap_8
XFILLER_111_602 VDD VSS sg13g2_decap_8
XFILLER_97_825 VDD VSS sg13g2_decap_8
X_2360_ _2360_/RESET_B VSS VDD _2360_/D _2360_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_110_112 VDD VSS sg13g2_decap_8
X_1311_ VDD _2185_/D _1311_/A VSS sg13g2_inv_1
XFILLER_2_770 VDD VSS sg13g2_decap_8
X_2291_ _2291_/RESET_B VSS VDD _2291_/D _2291_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_111_679 VDD VSS sg13g2_decap_8
XFILLER_96_357 VDD VSS sg13g2_decap_8
XFILLER_1_280 VDD VSS sg13g2_decap_8
XFILLER_2_42 VDD VSS sg13g2_decap_8
X_1242_ _1242_/B _2294_/Q _1249_/A VDD VSS sg13g2_xor2_1
XFILLER_77_593 VDD VSS sg13g2_decap_8
XFILLER_110_189 VDD VSS sg13g2_decap_8
XFILLER_38_947 VDD VSS sg13g2_decap_8
XFILLER_37_413 VDD VSS sg13g2_decap_8
XFILLER_65_766 VDD VSS sg13g2_decap_8
XFILLER_49_295 VDD VSS sg13g2_decap_8
XFILLER_80_725 VDD VSS sg13g2_decap_8
XFILLER_65_799 VDD VSS sg13g2_decap_8
XFILLER_64_254 VDD VSS sg13g2_decap_8
XFILLER_75_1010 VDD VSS sg13g2_decap_8
X_2271__213 VDD VSS _2271_/RESET_B sg13g2_tiehi
XFILLER_33_630 VDD VSS sg13g2_decap_8
XFILLER_52_438 VDD VSS sg13g2_decap_8
XFILLER_18_693 VDD VSS sg13g2_decap_8
XFILLER_45_490 VDD VSS sg13g2_decap_8
XFILLER_32_140 VDD VSS sg13g2_decap_8
XFILLER_21_847 VDD VSS sg13g2_decap_8
XFILLER_60_460 VDD VSS sg13g2_fill_1
XFILLER_20_357 VDD VSS sg13g2_decap_8
XFILLER_107_919 VDD VSS sg13g2_decap_8
XFILLER_106_407 VDD VSS sg13g2_decap_8
XFILLER_102_602 VDD VSS sg13g2_decap_8
XFILLER_99_151 VDD VSS sg13g2_fill_2
XFILLER_99_140 VDD VSS sg13g2_decap_8
XFILLER_0_707 VDD VSS sg13g2_decap_8
XFILLER_82_1047 VDD VSS sg13g2_decap_8
XFILLER_88_858 VDD VSS sg13g2_decap_8
XFILLER_99_184 VDD VSS sg13g2_decap_8
XFILLER_101_112 VDD VSS sg13g2_decap_8
X_1509_ _1671_/C _1509_/B _2270_/D VDD VSS sg13g2_nor2_1
XFILLER_29_903 VDD VSS sg13g2_decap_8
XFILLER_68_593 VDD VSS sg13g2_fill_2
XFILLER_56_700 VDD VSS sg13g2_decap_8
XFILLER_28_413 VDD VSS sg13g2_decap_8
XFILLER_110_690 VDD VSS sg13g2_decap_8
XFILLER_55_210 VDD VSS sg13g2_decap_8
XFILLER_83_585 VDD VSS sg13g2_decap_8
XFILLER_102_21 VDD VSS sg13g2_decap_8
XFILLER_44_928 VDD VSS sg13g2_decap_8
XFILLER_37_980 VDD VSS sg13g2_decap_8
XFILLER_56_777 VDD VSS sg13g2_decap_8
XFILLER_83_596 VDD VSS sg13g2_fill_1
XFILLER_24_630 VDD VSS sg13g2_decap_8
XFILLER_55_287 VDD VSS sg13g2_decap_8
XFILLER_36_490 VDD VSS sg13g2_decap_8
XFILLER_43_427 VDD VSS sg13g2_decap_8
XFILLER_52_950 VDD VSS sg13g2_fill_2
XFILLER_52_961 VDD VSS sg13g2_decap_4
XFILLER_23_140 VDD VSS sg13g2_decap_8
XFILLER_62_14 VDD VSS sg13g2_decap_8
XFILLER_102_98 VDD VSS sg13g2_decap_8
XFILLER_52_983 VDD VSS sg13g2_decap_8
XFILLER_12_847 VDD VSS sg13g2_decap_8
XFILLER_11_357 VDD VSS sg13g2_decap_8
XFILLER_109_212 VDD VSS sg13g2_fill_1
XFILLER_106_930 VDD VSS sg13g2_decap_8
XFILLER_11_84 VDD VSS sg13g2_decap_8
XFILLER_78_302 VDD VSS sg13g2_decap_8
XFILLER_3_567 VDD VSS sg13g2_decap_8
XFILLER_78_335 VDD VSS sg13g2_decap_8
XFILLER_78_313 VDD VSS sg13g2_fill_1
XFILLER_87_77 VDD VSS sg13g2_decap_8
XFILLER_78_368 VDD VSS sg13g2_decap_8
XFILLER_66_519 VDD VSS sg13g2_decap_8
XFILLER_59_560 VDD VSS sg13g2_decap_8
XFILLER_19_413 VDD VSS sg13g2_decap_8
XFILLER_98_1032 VDD VSS sg13g2_decap_8
XFILLER_4_1036 VDD VSS sg13g2_decap_8
XFILLER_74_574 VDD VSS sg13g2_decap_8
XFILLER_35_917 VDD VSS sg13g2_decap_8
XFILLER_28_980 VDD VSS sg13g2_decap_8
XFILLER_62_747 VDD VSS sg13g2_decap_8
XFILLER_61_213 VDD VSS sg13g2_decap_8
XFILLER_15_630 VDD VSS sg13g2_decap_8
XFILLER_36_70 VDD VSS sg13g2_decap_8
XFILLER_27_490 VDD VSS sg13g2_decap_8
XFILLER_34_427 VDD VSS sg13g2_decap_8
XFILLER_43_961 VDD VSS sg13g2_decap_8
XFILLER_61_246 VDD VSS sg13g2_decap_8
XFILLER_14_140 VDD VSS sg13g2_decap_8
XFILLER_70_780 VDD VSS sg13g2_decap_8
XFILLER_99_7 VDD VSS sg13g2_decap_8
X_1860_ _1860_/A _1907_/A _1952_/B VDD VSS sg13g2_and2_1
XFILLER_30_644 VDD VSS sg13g2_decap_8
X_1791_ _2223_/Q _2215_/Q _1812_/B VDD VSS sg13g2_xor2_1
XFILLER_7_840 VDD VSS sg13g2_decap_8
XFILLER_6_350 VDD VSS sg13g2_decap_8
XFILLER_69_302 VDD VSS sg13g2_decap_8
XFILLER_97_633 VDD VSS sg13g2_decap_8
X_2343_ _2343_/RESET_B VSS VDD _2343_/D _2343_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_112_966 VDD VSS sg13g2_decap_8
XFILLER_85_817 VDD VSS sg13g2_decap_8
XFILLER_96_154 VDD VSS sg13g2_decap_8
XFILLER_111_476 VDD VSS sg13g2_decap_8
XFILLER_69_379 VDD VSS sg13g2_decap_8
X_2274_ _2274_/RESET_B VSS VDD _2274_/D _2274_/Q _2289_/CLK sg13g2_dfrbpq_1
X_1225_ _1225_/X _2150_/A _1225_/B _2365_/Q VDD VSS sg13g2_and3_1
XFILLER_38_744 VDD VSS sg13g2_decap_8
XFILLER_37_210 VDD VSS sg13g2_decap_8
XFILLER_26_917 VDD VSS sg13g2_decap_8
XFILLER_53_725 VDD VSS sg13g2_decap_4
XFILLER_93_894 VDD VSS sg13g2_decap_8
XFILLER_80_544 VDD VSS sg13g2_decap_8
XFILLER_92_382 VDD VSS sg13g2_decap_8
XFILLER_19_980 VDD VSS sg13g2_decap_8
XFILLER_25_427 VDD VSS sg13g2_decap_8
XFILLER_37_287 VDD VSS sg13g2_decap_8
XFILLER_52_202 VDD VSS sg13g2_decap_8
XFILLER_80_577 VDD VSS sg13g2_decap_8
XFILLER_41_909 VDD VSS sg13g2_decap_8
XFILLER_18_490 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_17_clk clkbuf_leaf_0_clk/A clkload2/A VDD VSS sg13g2_buf_8
XFILLER_52_257 VDD VSS sg13g2_decap_4
XFILLER_34_994 VDD VSS sg13g2_decap_8
XFILLER_40_419 VDD VSS sg13g2_decap_8
XFILLER_21_644 VDD VSS sg13g2_decap_8
XFILLER_32_28 VDD VSS sg13g2_decap_8
XFILLER_20_154 VDD VSS sg13g2_decap_8
X_1989_ _2000_/C _2005_/B _2000_/B _1989_/Y VDD VSS sg13g2_nand3_1
XFILLER_107_716 VDD VSS sg13g2_decap_8
XFILLER_10_1008 VDD VSS sg13g2_decap_8
XFILLER_88_600 VDD VSS sg13g2_decap_8
XFILLER_106_259 VDD VSS sg13g2_decap_8
XFILLER_0_504 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[5\].out_data_pad out_data_PADs[5] bondpad_70x70
XFILLER_102_421 VDD VSS sg13g2_decap_8
XFILLER_102_410 VDD VSS sg13g2_decap_8
XFILLER_103_966 VDD VSS sg13g2_decap_8
XFILLER_57_14 VDD VSS sg13g2_decap_8
XFILLER_75_327 VDD VSS sg13g2_decap_8
XFILLER_87_165 VDD VSS sg13g2_decap_8
XFILLER_29_700 VDD VSS sg13g2_decap_8
XFILLER_102_498 VDD VSS sg13g2_decap_8
XFILLER_28_210 VDD VSS sg13g2_decap_8
XFILLER_90_319 VDD VSS sg13g2_decap_8
XFILLER_56_574 VDD VSS sg13g2_decap_8
XFILLER_29_777 VDD VSS sg13g2_decap_8
XFILLER_17_917 VDD VSS sg13g2_decap_8
X_2358__276 VDD VSS _2358_/RESET_B sg13g2_tiehi
XFILLER_73_35 VDD VSS sg13g2_decap_8
XFILLER_44_725 VDD VSS sg13g2_decap_8
XFILLER_16_427 VDD VSS sg13g2_decap_8
XFILLER_28_287 VDD VSS sg13g2_decap_8
XFILLER_43_224 VDD VSS sg13g2_decap_4
XFILLER_25_994 VDD VSS sg13g2_decap_8
XFILLER_19_1022 VDD VSS sg13g2_decap_8
XFILLER_43_279 VDD VSS sg13g2_fill_2
XFILLER_106_1014 VDD VSS sg13g2_decap_8
XFILLER_40_942 VDD VSS sg13g2_decap_8
XFILLER_12_644 VDD VSS sg13g2_decap_8
XFILLER_11_154 VDD VSS sg13g2_decap_8
XFILLER_8_637 VDD VSS sg13g2_decap_8
XFILLER_7_147 VDD VSS sg13g2_decap_8
XFILLER_98_21 VDD VSS sg13g2_decap_8
X_2365__269 VDD VSS _2365_/RESET_B sg13g2_tiehi
XFILLER_4_854 VDD VSS sg13g2_decap_8
XFILLER_105_270 VDD VSS sg13g2_decap_8
XFILLER_98_98 VDD VSS sg13g2_decap_8
XFILLER_3_364 VDD VSS sg13g2_decap_8
XFILLER_105_281 VDD VSS sg13g2_fill_1
XFILLER_26_1015 VDD VSS sg13g2_decap_8
XFILLER_94_636 VDD VSS sg13g2_decap_4
XFILLER_79_699 VDD VSS sg13g2_decap_4
XFILLER_78_154 VDD VSS sg13g2_decap_4
XFILLER_94_669 VDD VSS sg13g2_decap_8
XFILLER_59_390 VDD VSS sg13g2_decap_8
XFILLER_14_7 VDD VSS sg13g2_decap_8
XFILLER_19_210 VDD VSS sg13g2_decap_8
XFILLER_75_883 VDD VSS sg13g2_decap_8
XFILLER_81_319 VDD VSS sg13g2_decap_8
XFILLER_47_552 VDD VSS sg13g2_fill_2
XFILLER_35_714 VDD VSS sg13g2_decap_8
XFILLER_62_500 VDD VSS sg13g2_fill_1
XFILLER_47_91 VDD VSS sg13g2_decap_8
XFILLER_90_820 VDD VSS sg13g2_decap_8
XFILLER_74_382 VDD VSS sg13g2_decap_8
XFILLER_62_533 VDD VSS sg13g2_decap_8
XFILLER_62_511 VDD VSS sg13g2_fill_1
XFILLER_19_287 VDD VSS sg13g2_decap_8
XFILLER_34_224 VDD VSS sg13g2_decap_8
XFILLER_16_994 VDD VSS sg13g2_decap_8
XFILLER_72_1046 VDD VSS sg13g2_decap_8
X_1912_ _1914_/A _1912_/A _1912_/B VDD VSS sg13g2_xnor2_1
XFILLER_33_1008 VDD VSS sg13g2_decap_8
XFILLER_31_931 VDD VSS sg13g2_decap_8
XFILLER_63_90 VDD VSS sg13g2_decap_8
XFILLER_30_441 VDD VSS sg13g2_decap_8
X_1843_ _1934_/B _1934_/A _1839_/Y _1843_/X VDD VSS sg13g2_a21o_1
XFILLER_8_63 VDD VSS sg13g2_decap_8
X_1774_ _1774_/B _1774_/A _1775_/B VDD VSS sg13g2_xor2_1
Xclkbuf_leaf_6_clk clkbuf_leaf_9_clk/A _2372_/CLK VDD VSS sg13g2_buf_8
XFILLER_103_207 VDD VSS sg13g2_fill_1
XFILLER_89_419 VDD VSS sg13g2_decap_8
XFILLER_98_931 VDD VSS sg13g2_decap_8
XFILLER_40_0 VDD VSS sg13g2_decap_8
XFILLER_112_763 VDD VSS sg13g2_decap_8
XFILLER_97_452 VDD VSS sg13g2_decap_8
XFILLER_98_997 VDD VSS sg13g2_fill_2
XFILLER_85_603 VDD VSS sg13g2_decap_8
X_2326_ _2326_/RESET_B VSS VDD _2326_/D _2326_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_111_273 VDD VSS sg13g2_decap_8
XFILLER_57_316 VDD VSS sg13g2_decap_8
XFILLER_84_135 VDD VSS sg13g2_decap_8
X_2257_ _2257_/RESET_B VSS VDD _2257_/D _2257_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_26_714 VDD VSS sg13g2_decap_8
X_1208_ VDD _1208_/Y _2210_/Q VSS sg13g2_inv_1
XFILLER_27_28 VDD VSS sg13g2_decap_8
XFILLER_81_842 VDD VSS sg13g2_decap_8
X_2188_ _2188_/RESET_B VSS VDD _2188_/D _2188_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_65_371 VDD VSS sg13g2_decap_8
XFILLER_25_224 VDD VSS sg13g2_decap_8
XFILLER_80_341 VDD VSS sg13g2_decap_8
XFILLER_53_566 VDD VSS sg13g2_decap_8
XFILLER_41_706 VDD VSS sg13g2_decap_8
XFILLER_22_931 VDD VSS sg13g2_decap_8
XFILLER_34_791 VDD VSS sg13g2_decap_8
XFILLER_43_49 VDD VSS sg13g2_decap_8
XFILLER_21_441 VDD VSS sg13g2_decap_8
XFILLER_108_42 VDD VSS sg13g2_decap_8
XFILLER_0_301 VDD VSS sg13g2_decap_8
XFILLER_68_35 VDD VSS sg13g2_decap_8
XFILLER_1_868 VDD VSS sg13g2_decap_8
XFILLER_76_603 VDD VSS sg13g2_decap_8
XFILLER_88_485 VDD VSS sg13g2_decap_8
XFILLER_49_839 VDD VSS sg13g2_decap_4
XFILLER_0_378 VDD VSS sg13g2_decap_8
XFILLER_88_496 VDD VSS sg13g2_fill_2
XFILLER_64_809 VDD VSS sg13g2_decap_8
XFILLER_84_56 VDD VSS sg13g2_decap_8
XFILLER_57_850 VDD VSS sg13g2_fill_2
XFILLER_17_714 VDD VSS sg13g2_decap_8
XFILLER_72_842 VDD VSS sg13g2_decap_8
XFILLER_90_105 VDD VSS sg13g2_decap_8
XFILLER_57_894 VDD VSS sg13g2_decap_8
XFILLER_29_574 VDD VSS sg13g2_decap_8
XFILLER_16_224 VDD VSS sg13g2_decap_8
XFILLER_44_522 VDD VSS sg13g2_decap_8
XFILLER_95_1057 VDD VSS sg13g2_decap_4
XFILLER_71_385 VDD VSS sg13g2_decap_8
XFILLER_44_599 VDD VSS sg13g2_decap_8
XFILLER_32_728 VDD VSS sg13g2_decap_8
XFILLER_25_791 VDD VSS sg13g2_decap_8
XFILLER_13_931 VDD VSS sg13g2_decap_8
XFILLER_31_238 VDD VSS sg13g2_decap_8
XFILLER_12_441 VDD VSS sg13g2_decap_8
XFILLER_9_924 VDD VSS sg13g2_decap_8
XFILLER_8_434 VDD VSS sg13g2_decap_8
XFILLER_4_651 VDD VSS sg13g2_decap_8
X_1490_ VSS VDD _1365_/B _2355_/Q _1490_/Y hold555/X sg13g2_a21oi_1
XFILLER_3_161 VDD VSS sg13g2_decap_8
XFILLER_67_614 VDD VSS sg13g2_decap_8
XFILLER_95_945 VDD VSS sg13g2_decap_8
XFILLER_94_433 VDD VSS sg13g2_decap_8
X_2111_ hold530/X VDD _2111_/Y VSS _1510_/A hold379/X sg13g2_o21ai_1
XFILLER_66_135 VDD VSS sg13g2_fill_1
XFILLER_39_338 VDD VSS sg13g2_decap_8
X_2042_ _2040_/Y VDD _2327_/D VSS _2156_/A _2041_/Y sg13g2_o21ai_1
XFILLER_66_146 VDD VSS sg13g2_decap_8
XFILLER_82_639 VDD VSS sg13g2_decap_8
XFILLER_81_105 VDD VSS sg13g2_decap_8
XFILLER_35_511 VDD VSS sg13g2_decap_8
XFILLER_47_371 VDD VSS sg13g2_decap_8
XFILLER_63_853 VDD VSS sg13g2_decap_8
XFILLER_62_330 VDD VSS sg13g2_decap_8
XFILLER_90_661 VDD VSS sg13g2_decap_8
XFILLER_35_588 VDD VSS sg13g2_decap_8
XFILLER_23_728 VDD VSS sg13g2_decap_8
XFILLER_50_525 VDD VSS sg13g2_decap_8
XFILLER_16_791 VDD VSS sg13g2_decap_8
XFILLER_22_238 VDD VSS sg13g2_decap_8
XFILLER_88_0 VDD VSS sg13g2_decap_8
X_1826_ _1826_/B _1826_/A _1827_/A VDD VSS sg13g2_xor2_1
Xhold401 _2197_/Q VDD VSS hold401/X sg13g2_dlygate4sd3_1
Xhold434 _1654_/Y VDD VSS _1655_/B sg13g2_dlygate4sd3_1
X_1757_ _1761_/B _1751_/X _1749_/A _1772_/B VDD VSS sg13g2_a21o_1
XFILLER_104_505 VDD VSS sg13g2_decap_4
Xhold412 _2227_/Q VDD VSS _1412_/A sg13g2_dlygate4sd3_1
Xhold445 _2247_/Q VDD VSS _1455_/A sg13g2_dlygate4sd3_1
Xhold423 _1669_/Y VDD VSS _1670_/B sg13g2_dlygate4sd3_1
Xhold467 _1700_/Y VDD VSS _1701_/B sg13g2_dlygate4sd3_1
XFILLER_104_538 VDD VSS sg13g2_decap_8
Xhold456 _2223_/Q VDD VSS hold456/X sg13g2_dlygate4sd3_1
X_1688_ _1725_/A _1688_/B _2307_/Q VDD VSS sg13g2_nand2b_1
Xhold478 _2278_/Q VDD VSS hold478/X sg13g2_dlygate4sd3_1
XFILLER_104_549 VDD VSS sg13g2_decap_8
Xhold489 _2234_/Q VDD VSS _1426_/A sg13g2_dlygate4sd3_1
XFILLER_86_923 VDD VSS sg13g2_decap_8
XFILLER_112_560 VDD VSS sg13g2_decap_8
XFILLER_98_794 VDD VSS sg13g2_fill_1
XFILLER_85_411 VDD VSS sg13g2_fill_2
XFILLER_58_658 VDD VSS sg13g2_decap_8
X_2309_ _2309__79/L_HI VSS VDD _2309_/D _2309_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_38_49 VDD VSS sg13g2_decap_8
XFILLER_86_989 VDD VSS sg13g2_decap_8
XFILLER_79_1008 VDD VSS sg13g2_decap_8
XFILLER_39_850 VDD VSS sg13g2_decap_8
XFILLER_57_157 VDD VSS sg13g2_decap_8
XFILLER_45_308 VDD VSS sg13g2_decap_8
XFILLER_73_639 VDD VSS sg13g2_decap_8
XFILLER_57_179 VDD VSS sg13g2_decap_8
XFILLER_26_511 VDD VSS sg13g2_decap_8
XFILLER_54_864 VDD VSS sg13g2_decap_8
XFILLER_26_588 VDD VSS sg13g2_decap_8
XFILLER_14_728 VDD VSS sg13g2_decap_8
XFILLER_0_1050 VDD VSS sg13g2_decap_8
XFILLER_54_59 VDD VSS sg13g2_fill_1
XFILLER_41_525 VDD VSS sg13g2_fill_1
XFILLER_81_694 VDD VSS sg13g2_decap_8
XFILLER_80_171 VDD VSS sg13g2_decap_8
XFILLER_110_21 VDD VSS sg13g2_decap_8
XFILLER_53_396 VDD VSS sg13g2_decap_8
XFILLER_13_238 VDD VSS sg13g2_decap_8
XFILLER_70_14 VDD VSS sg13g2_decap_8
XFILLER_55_1052 VDD VSS sg13g2_decap_8
XFILLER_110_98 VDD VSS sg13g2_decap_8
XFILLER_10_945 VDD VSS sg13g2_decap_8
XFILLER_16_1036 VDD VSS sg13g2_decap_8
XFILLER_108_822 VDD VSS sg13g2_decap_8
XFILLER_6_938 VDD VSS sg13g2_decap_8
XFILLER_107_332 VDD VSS sg13g2_decap_8
XFILLER_5_448 VDD VSS sg13g2_decap_8
XFILLER_108_899 VDD VSS sg13g2_decap_8
XFILLER_79_56 VDD VSS sg13g2_decap_8
XFILLER_77_912 VDD VSS sg13g2_decap_8
XFILLER_110_508 VDD VSS sg13g2_decap_8
XFILLER_1_665 VDD VSS sg13g2_decap_8
XFILLER_76_422 VDD VSS sg13g2_decap_8
XFILLER_23_1029 VDD VSS sg13g2_decap_8
XFILLER_49_636 VDD VSS sg13g2_fill_2
XFILLER_0_175 VDD VSS sg13g2_decap_8
XFILLER_91_403 VDD VSS sg13g2_decap_8
XFILLER_76_455 VDD VSS sg13g2_decap_8
XFILLER_95_77 VDD VSS sg13g2_decap_8
XFILLER_64_606 VDD VSS sg13g2_decap_8
XFILLER_48_146 VDD VSS sg13g2_decap_4
XFILLER_36_308 VDD VSS sg13g2_decap_8
XFILLER_48_168 VDD VSS sg13g2_decap_8
XFILLER_91_414 VDD VSS sg13g2_fill_2
XFILLER_17_511 VDD VSS sg13g2_decap_8
XFILLER_63_127 VDD VSS sg13g2_fill_1
XFILLER_29_371 VDD VSS sg13g2_decap_8
XFILLER_91_447 VDD VSS sg13g2_decap_8
XFILLER_63_138 VDD VSS sg13g2_decap_8
X_2217__106 VDD VSS _2217_/RESET_B sg13g2_tiehi
XFILLER_17_588 VDD VSS sg13g2_decap_8
XFILLER_60_834 VDD VSS sg13g2_fill_1
XFILLER_44_70 VDD VSS sg13g2_decap_8
XFILLER_32_525 VDD VSS sg13g2_decap_8
XFILLER_44_385 VDD VSS sg13g2_decap_8
XFILLER_81_7 VDD VSS sg13g2_decap_8
XFILLER_9_721 VDD VSS sg13g2_decap_8
XFILLER_8_231 VDD VSS sg13g2_decap_8
XFILLER_9_798 VDD VSS sg13g2_decap_8
X_1611_ _1617_/A _2292_/Q _2277_/Q VDD VSS sg13g2_xnor2_1
XFILLER_60_80 VDD VSS sg13g2_decap_8
X_1542_ _1556_/S0 _2237_/Q _2229_/Q _2221_/Q _2213_/Q _1589_/B _1543_/A VDD VSS sg13g2_mux4_1
XFILLER_5_42 VDD VSS sg13g2_decap_8
XFILLER_99_569 VDD VSS sg13g2_decap_8
X_1473_ VSS VDD _1198_/Y _1465_/Y _1473_/Y _1472_/Y sg13g2_a21oi_1
X_2163__271 VDD VSS _2163_/RESET_B sg13g2_tiehi
XFILLER_67_422 VDD VSS sg13g2_decap_8
XFILLER_27_308 VDD VSS sg13g2_decap_8
XFILLER_39_168 VDD VSS sg13g2_decap_8
XFILLER_94_296 VDD VSS sg13g2_decap_8
XFILLER_82_436 VDD VSS sg13g2_decap_8
XFILLER_48_680 VDD VSS sg13g2_decap_8
XFILLER_54_127 VDD VSS sg13g2_decap_8
X_2025_ _2025_/A _2024_/X _2025_/Y VDD VSS sg13g2_nor2b_1
XFILLER_39_1025 VDD VSS sg13g2_decap_8
XFILLER_36_875 VDD VSS sg13g2_decap_8
XFILLER_23_525 VDD VSS sg13g2_decap_8
XFILLER_35_385 VDD VSS sg13g2_decap_8
XFILLER_50_311 VDD VSS sg13g2_decap_8
XFILLER_51_867 VDD VSS sg13g2_decap_8
XFILLER_51_878 VDD VSS sg13g2_fill_1
XFILLER_50_388 VDD VSS sg13g2_decap_8
XFILLER_40_28 VDD VSS sg13g2_decap_8
XFILLER_85_1001 VDD VSS sg13g2_fill_2
X_1809_ _1930_/A _1809_/A _1809_/B VDD VSS sg13g2_nand2_1
XFILLER_85_1023 VDD VSS sg13g2_fill_2
XFILLER_105_847 VDD VSS sg13g2_decap_8
XFILLER_104_335 VDD VSS sg13g2_decap_8
XFILLER_59_901 VDD VSS sg13g2_decap_8
Xhold297 _2285_/Q VDD VSS _1226_/B sg13g2_dlygate4sd3_1
XFILLER_105_21 VDD VSS sg13g2_decap_8
XFILLER_74_926 VDD VSS sg13g2_decap_8
XFILLER_86_753 VDD VSS sg13g2_decap_8
XFILLER_85_252 VDD VSS sg13g2_decap_8
XFILLER_59_978 VDD VSS sg13g2_decap_8
XFILLER_18_308 VDD VSS sg13g2_decap_8
XFILLER_65_14 VDD VSS sg13g2_decap_8
XFILLER_100_574 VDD VSS sg13g2_decap_8
XFILLER_73_414 VDD VSS sg13g2_decap_8
XFILLER_105_98 VDD VSS sg13g2_decap_8
XFILLER_46_628 VDD VSS sg13g2_fill_1
XFILLER_82_970 VDD VSS sg13g2_decap_8
XFILLER_82_981 VDD VSS sg13g2_fill_2
XFILLER_54_661 VDD VSS sg13g2_decap_8
XFILLER_42_812 VDD VSS sg13g2_decap_8
XFILLER_27_875 VDD VSS sg13g2_decap_8
XFILLER_92_1049 VDD VSS sg13g2_decap_8
XFILLER_92_1038 VDD VSS sg13g2_fill_2
XFILLER_81_35 VDD VSS sg13g2_decap_8
XFILLER_53_182 VDD VSS sg13g2_decap_8
XFILLER_14_525 VDD VSS sg13g2_decap_8
XFILLER_26_385 VDD VSS sg13g2_decap_8
XFILLER_41_322 VDD VSS sg13g2_decap_8
XFILLER_42_889 VDD VSS sg13g2_decap_8
XFILLER_41_388 VDD VSS sg13g2_decap_8
XFILLER_14_84 VDD VSS sg13g2_decap_8
XFILLER_10_742 VDD VSS sg13g2_decap_8
XFILLER_6_735 VDD VSS sg13g2_decap_8
XFILLER_5_245 VDD VSS sg13g2_decap_8
XFILLER_108_696 VDD VSS sg13g2_decap_8
XFILLER_107_140 VDD VSS sg13g2_decap_8
XFILLER_2_952 VDD VSS sg13g2_decap_8
XFILLER_96_528 VDD VSS sg13g2_decap_8
XFILLER_1_462 VDD VSS sg13g2_decap_8
XFILLER_7_1001 VDD VSS sg13g2_decap_8
XFILLER_49_433 VDD VSS sg13g2_decap_8
XFILLER_77_753 VDD VSS sg13g2_decap_8
XFILLER_103_390 VDD VSS sg13g2_decap_8
XFILLER_39_70 VDD VSS sg13g2_decap_8
XFILLER_65_937 VDD VSS sg13g2_decap_8
XFILLER_36_105 VDD VSS sg13g2_decap_8
XFILLER_92_756 VDD VSS sg13g2_decap_8
XFILLER_76_296 VDD VSS sg13g2_fill_2
XFILLER_64_458 VDD VSS sg13g2_decap_8
XFILLER_91_255 VDD VSS sg13g2_decap_8
XFILLER_33_812 VDD VSS sg13g2_decap_8
XFILLER_18_875 VDD VSS sg13g2_decap_8
XFILLER_51_119 VDD VSS sg13g2_decap_8
XFILLER_45_683 VDD VSS sg13g2_decap_8
XFILLER_17_385 VDD VSS sg13g2_decap_8
XFILLER_32_322 VDD VSS sg13g2_decap_8
XFILLER_33_889 VDD VSS sg13g2_decap_8
XFILLER_44_193 VDD VSS sg13g2_decap_8
XFILLER_60_686 VDD VSS sg13g2_fill_2
XFILLER_20_539 VDD VSS sg13g2_decap_8
XFILLER_32_399 VDD VSS sg13g2_decap_8
XFILLER_9_595 VDD VSS sg13g2_decap_8
XFILLER_99_311 VDD VSS sg13g2_decap_8
X_1525_ _1527_/B _1576_/A _2284_/D VDD VSS sg13g2_nor2_1
XFILLER_102_806 VDD VSS sg13g2_fill_1
XFILLER_59_208 VDD VSS sg13g2_decap_8
XFILLER_102_839 VDD VSS sg13g2_decap_8
XFILLER_101_316 VDD VSS sg13g2_decap_8
X_1456_ VSS VDD _1376_/Y _1455_/B _2247_/D _1455_/Y sg13g2_a21oi_1
XFILLER_95_561 VDD VSS sg13g2_decap_8
X_1387_ _1386_/Y VDD _2217_/D VSS _1367_/B _1385_/Y sg13g2_o21ai_1
XFILLER_68_764 VDD VSS sg13g2_decap_8
XFILLER_67_230 VDD VSS sg13g2_decap_8
XFILLER_110_872 VDD VSS sg13g2_decap_8
XFILLER_83_712 VDD VSS sg13g2_decap_8
XFILLER_56_948 VDD VSS sg13g2_fill_2
XFILLER_27_105 VDD VSS sg13g2_decap_8
XFILLER_71_907 VDD VSS sg13g2_decap_8
XFILLER_82_222 VDD VSS sg13g2_decap_8
XFILLER_36_672 VDD VSS sg13g2_decap_8
XFILLER_24_812 VDD VSS sg13g2_decap_8
XFILLER_35_28 VDD VSS sg13g2_decap_8
X_2008_ _1931_/A _1901_/B _2021_/S _2008_/X VDD VSS sg13g2_mux2_1
XFILLER_82_299 VDD VSS sg13g2_decap_8
XFILLER_42_119 VDD VSS sg13g2_decap_8
XFILLER_23_322 VDD VSS sg13g2_decap_8
XFILLER_35_182 VDD VSS sg13g2_decap_8
XFILLER_51_675 VDD VSS sg13g2_decap_8
XFILLER_24_889 VDD VSS sg13g2_decap_8
XFILLER_91_1060 VDD VSS sg13g2_fill_1
XFILLER_52_1011 VDD VSS sg13g2_decap_8
XFILLER_52_1022 VDD VSS sg13g2_fill_2
XFILLER_11_539 VDD VSS sg13g2_decap_8
XFILLER_23_399 VDD VSS sg13g2_decap_8
XFILLER_50_174 VDD VSS sg13g2_decap_8
XFILLER_109_427 VDD VSS sg13g2_decap_8
Xout_data_pads\[2\].out_data_pad _2368_/Q IOVDD IOVSS out_data_PADs[2] VDD VSS sg13g2_IOPadOut30mA
XFILLER_105_644 VDD VSS sg13g2_decap_8
XFILLER_3_749 VDD VSS sg13g2_decap_8
XFILLER_2_259 VDD VSS sg13g2_decap_8
XFILLER_76_35 VDD VSS sg13g2_decap_8
XFILLER_59_742 VDD VSS sg13g2_decap_8
XFILLER_47_915 VDD VSS sg13g2_decap_8
XFILLER_58_241 VDD VSS sg13g2_decap_8
XFILLER_101_883 VDD VSS sg13g2_decap_8
XFILLER_58_252 VDD VSS sg13g2_fill_2
XFILLER_18_105 VDD VSS sg13g2_decap_8
XFILLER_46_414 VDD VSS sg13g2_fill_2
XFILLER_73_222 VDD VSS sg13g2_decap_8
XFILLER_73_277 VDD VSS sg13g2_decap_4
XFILLER_34_609 VDD VSS sg13g2_decap_8
XFILLER_27_672 VDD VSS sg13g2_decap_8
XFILLER_15_812 VDD VSS sg13g2_decap_8
X_2292__141 VDD VSS _2292_/RESET_B sg13g2_tiehi
XFILLER_109_1001 VDD VSS sg13g2_decap_8
XFILLER_73_299 VDD VSS sg13g2_fill_1
XFILLER_92_56 VDD VSS sg13g2_decap_8
XFILLER_61_439 VDD VSS sg13g2_decap_8
XFILLER_14_322 VDD VSS sg13g2_decap_8
XFILLER_33_119 VDD VSS sg13g2_decap_8
XFILLER_26_182 VDD VSS sg13g2_decap_8
XFILLER_70_962 VDD VSS sg13g2_decap_8
XFILLER_15_889 VDD VSS sg13g2_decap_8
XFILLER_42_686 VDD VSS sg13g2_decap_8
XFILLER_30_826 VDD VSS sg13g2_decap_8
XFILLER_14_399 VDD VSS sg13g2_decap_8
XFILLER_41_174 VDD VSS sg13g2_decap_8
XFILLER_6_532 VDD VSS sg13g2_decap_8
XFILLER_109_994 VDD VSS sg13g2_decap_8
XFILLER_108_471 VDD VSS sg13g2_decap_8
XFILLER_68_1040 VDD VSS sg13g2_decap_8
XFILLER_44_7 VDD VSS sg13g2_decap_8
XFILLER_29_1057 VDD VSS sg13g2_decap_4
XFILLER_96_336 VDD VSS sg13g2_decap_8
X_1310_ _1310_/Y _1482_/B1 hold383/X _1482_/A2 _2349_/Q VDD VSS sg13g2_a22oi_1
X_2290_ _2290_/RESET_B VSS VDD _2290_/D _2290_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_111_658 VDD VSS sg13g2_decap_8
XFILLER_2_21 VDD VSS sg13g2_decap_8
X_1241_ _1247_/A _2293_/Q _2255_/Q VDD VSS sg13g2_xnor2_1
XFILLER_77_572 VDD VSS sg13g2_decap_8
XFILLER_110_168 VDD VSS sg13g2_decap_8
XFILLER_38_926 VDD VSS sg13g2_decap_8
XFILLER_49_274 VDD VSS sg13g2_decap_8
XFILLER_65_745 VDD VSS sg13g2_decap_8
XFILLER_64_233 VDD VSS sg13g2_decap_8
XFILLER_2_98 VDD VSS sg13g2_decap_8
XFILLER_92_586 VDD VSS sg13g2_decap_8
XFILLER_53_918 VDD VSS sg13g2_decap_8
XFILLER_25_609 VDD VSS sg13g2_decap_8
XFILLER_52_417 VDD VSS sg13g2_fill_2
XFILLER_18_672 VDD VSS sg13g2_decap_8
XFILLER_37_469 VDD VSS sg13g2_decap_8
XFILLER_17_182 VDD VSS sg13g2_decap_8
XFILLER_24_119 VDD VSS sg13g2_decap_8
XFILLER_61_951 VDD VSS sg13g2_decap_8
XFILLER_61_995 VDD VSS sg13g2_fill_1
XFILLER_33_686 VDD VSS sg13g2_decap_8
XFILLER_21_826 VDD VSS sg13g2_decap_8
XFILLER_20_336 VDD VSS sg13g2_decap_8
XFILLER_32_196 VDD VSS sg13g2_decap_8
XFILLER_70_0 VDD VSS sg13g2_decap_8
XFILLER_9_392 VDD VSS sg13g2_decap_8
XFILLER_12_1050 VDD VSS sg13g2_decap_8
XFILLER_82_1026 VDD VSS sg13g2_decap_8
XFILLER_99_163 VDD VSS sg13g2_decap_8
XFILLER_88_837 VDD VSS sg13g2_decap_8
X_1508_ _1509_/B _1506_/X _1507_/Y _1503_/X _1510_/B VDD VSS sg13g2_a22oi_1
X_1439_ VDD _2239_/D _1439_/A VSS sg13g2_inv_1
XFILLER_96_892 VDD VSS sg13g2_decap_8
XFILLER_101_179 VDD VSS sg13g2_decap_4
XFILLER_68_572 VDD VSS sg13g2_decap_8
XFILLER_83_520 VDD VSS sg13g2_fill_1
XFILLER_29_959 VDD VSS sg13g2_decap_8
XFILLER_56_756 VDD VSS sg13g2_decap_8
XFILLER_44_907 VDD VSS sg13g2_decap_8
XFILLER_46_49 VDD VSS sg13g2_decap_8
XFILLER_83_564 VDD VSS sg13g2_decap_8
XFILLER_55_266 VDD VSS sg13g2_decap_8
XFILLER_16_609 VDD VSS sg13g2_decap_8
XFILLER_28_469 VDD VSS sg13g2_decap_8
XFILLER_43_406 VDD VSS sg13g2_decap_8
XFILLER_71_748 VDD VSS sg13g2_decap_8
XFILLER_70_236 VDD VSS sg13g2_fill_2
XFILLER_15_119 VDD VSS sg13g2_decap_8
XFILLER_102_77 VDD VSS sg13g2_decap_8
XFILLER_24_686 VDD VSS sg13g2_decap_8
XFILLER_51_483 VDD VSS sg13g2_decap_8
XFILLER_51_450 VDD VSS sg13g2_fill_1
XFILLER_12_826 VDD VSS sg13g2_decap_8
XFILLER_51_494 VDD VSS sg13g2_fill_2
XFILLER_11_336 VDD VSS sg13g2_decap_8
XFILLER_8_819 VDD VSS sg13g2_decap_8
XFILLER_23_196 VDD VSS sg13g2_decap_8
XFILLER_7_329 VDD VSS sg13g2_decap_8
XFILLER_109_279 VDD VSS sg13g2_decap_8
XFILLER_11_63 VDD VSS sg13g2_decap_8
XFILLER_3_546 VDD VSS sg13g2_decap_8
XFILLER_106_986 VDD VSS sg13g2_decap_8
XFILLER_105_463 VDD VSS sg13g2_decap_8
XFILLER_87_56 VDD VSS sg13g2_decap_8
XFILLER_94_829 VDD VSS sg13g2_decap_8
XFILLER_93_317 VDD VSS sg13g2_decap_8
XFILLER_47_712 VDD VSS sg13g2_decap_8
XFILLER_4_1015 VDD VSS sg13g2_decap_8
XFILLER_86_391 VDD VSS sg13g2_decap_8
XFILLER_74_553 VDD VSS sg13g2_decap_8
XFILLER_59_1028 VDD VSS sg13g2_fill_2
XFILLER_59_1006 VDD VSS sg13g2_decap_8
XFILLER_47_778 VDD VSS sg13g2_decap_4
XFILLER_19_469 VDD VSS sg13g2_decap_8
XFILLER_34_406 VDD VSS sg13g2_decap_8
XFILLER_62_726 VDD VSS sg13g2_decap_8
XFILLER_46_277 VDD VSS sg13g2_decap_8
XFILLER_43_940 VDD VSS sg13g2_decap_8
XFILLER_30_623 VDD VSS sg13g2_decap_8
XFILLER_15_686 VDD VSS sg13g2_decap_8
XFILLER_42_461 VDD VSS sg13g2_decap_8
XFILLER_35_1050 VDD VSS sg13g2_decap_8
XFILLER_14_196 VDD VSS sg13g2_decap_8
X_1790_ _1801_/A _2223_/Q _2215_/Q VDD VSS sg13g2_nand2b_1
XIO_FILL_IO_WEST_1_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_109_791 VDD VSS sg13g2_decap_8
XFILLER_7_896 VDD VSS sg13g2_decap_8
XFILLER_112_945 VDD VSS sg13g2_decap_8
X_2342_ _2342_/RESET_B VSS VDD _2342_/D _2342_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_111_455 VDD VSS sg13g2_decap_8
XFILLER_96_133 VDD VSS sg13g2_decap_8
XFILLER_78_881 VDD VSS sg13g2_decap_8
XFILLER_84_306 VDD VSS sg13g2_decap_8
XFILLER_42_1043 VDD VSS sg13g2_decap_8
X_2273_ _2273_/RESET_B VSS VDD _2273_/D _2273_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_38_723 VDD VSS sg13g2_decap_8
XFILLER_77_391 VDD VSS sg13g2_decap_8
X_1224_ _2150_/A _1502_/D _2360_/D VDD VSS sg13g2_and2_1
XFILLER_93_873 VDD VSS sg13g2_decap_8
XFILLER_93_884 VDD VSS sg13g2_fill_1
XFILLER_92_361 VDD VSS sg13g2_decap_8
XFILLER_65_564 VDD VSS sg13g2_decap_8
XFILLER_53_704 VDD VSS sg13g2_decap_8
XFILLER_25_406 VDD VSS sg13g2_decap_8
XFILLER_37_266 VDD VSS sg13g2_decap_8
XFILLER_80_523 VDD VSS sg13g2_decap_8
XFILLER_52_236 VDD VSS sg13g2_decap_8
XFILLER_34_973 VDD VSS sg13g2_decap_8
XFILLER_21_623 VDD VSS sg13g2_decap_8
XFILLER_60_291 VDD VSS sg13g2_decap_4
XFILLER_33_483 VDD VSS sg13g2_decap_8
XFILLER_20_133 VDD VSS sg13g2_decap_8
X_1988_ _2005_/B _1988_/A _1988_/B VDD VSS sg13g2_nand2_1
XFILLER_106_238 VDD VSS sg13g2_decap_8
XFILLER_103_945 VDD VSS sg13g2_decap_8
XFILLER_87_144 VDD VSS sg13g2_decap_8
XFILLER_102_477 VDD VSS sg13g2_decap_8
XFILLER_75_306 VDD VSS sg13g2_decap_8
XFILLER_29_756 VDD VSS sg13g2_decap_8
Xclkbuf_2_2__f_clk clkbuf_2_2__f_clk/X clkbuf_0_clk/X VDD VSS sg13g2_buf_16
XFILLER_44_704 VDD VSS sg13g2_decap_8
XFILLER_16_406 VDD VSS sg13g2_decap_8
XFILLER_28_266 VDD VSS sg13g2_decap_8
XFILLER_73_14 VDD VSS sg13g2_decap_8
XFILLER_43_203 VDD VSS sg13g2_decap_8
XFILLER_19_1001 VDD VSS sg13g2_decap_8
XFILLER_43_258 VDD VSS sg13g2_decap_8
XFILLER_40_921 VDD VSS sg13g2_decap_8
XFILLER_25_973 VDD VSS sg13g2_decap_8
XFILLER_12_623 VDD VSS sg13g2_decap_8
XFILLER_24_483 VDD VSS sg13g2_decap_8
XFILLER_40_998 VDD VSS sg13g2_decap_8
XFILLER_11_133 VDD VSS sg13g2_decap_8
XFILLER_8_616 VDD VSS sg13g2_decap_8
XFILLER_7_126 VDD VSS sg13g2_decap_8
XFILLER_22_84 VDD VSS sg13g2_decap_8
XFILLER_4_833 VDD VSS sg13g2_decap_8
XFILLER_98_77 VDD VSS sg13g2_decap_8
XFILLER_3_343 VDD VSS sg13g2_decap_8
XFILLER_106_783 VDD VSS sg13g2_decap_8
XFILLER_65_1043 VDD VSS sg13g2_decap_8
XFILLER_0_0 VDD VSS sg13g2_decap_8
XFILLER_78_133 VDD VSS sg13g2_decap_8
XFILLER_94_615 VDD VSS sg13g2_decap_8
XFILLER_79_678 VDD VSS sg13g2_decap_8
XFILLER_78_199 VDD VSS sg13g2_decap_8
XFILLER_75_862 VDD VSS sg13g2_decap_8
XFILLER_93_147 VDD VSS sg13g2_decap_8
XFILLER_47_564 VDD VSS sg13g2_decap_8
XFILLER_47_597 VDD VSS sg13g2_fill_1
XFILLER_19_266 VDD VSS sg13g2_decap_8
XFILLER_34_203 VDD VSS sg13g2_decap_8
XFILLER_90_865 VDD VSS sg13g2_decap_8
XFILLER_50_718 VDD VSS sg13g2_decap_8
XFILLER_31_910 VDD VSS sg13g2_decap_8
XFILLER_16_973 VDD VSS sg13g2_decap_8
XFILLER_72_1025 VDD VSS sg13g2_decap_8
X_1911_ VSS VDD _1985_/A _1911_/B _1911_/A sg13g2_or2_1
XFILLER_15_483 VDD VSS sg13g2_decap_8
XFILLER_30_420 VDD VSS sg13g2_decap_8
XFILLER_42_280 VDD VSS sg13g2_decap_8
X_1842_ VSS VDD _1934_/A _1934_/B _1905_/B _1839_/Y sg13g2_a21oi_1
XFILLER_31_987 VDD VSS sg13g2_decap_8
XFILLER_8_42 VDD VSS sg13g2_decap_8
XFILLER_30_497 VDD VSS sg13g2_decap_8
X_1773_ _1877_/A VDD _1775_/A VSS _1927_/A _1877_/B sg13g2_o21ai_1
XFILLER_7_693 VDD VSS sg13g2_decap_8
XFILLER_98_976 VDD VSS sg13g2_decap_8
XFILLER_112_742 VDD VSS sg13g2_decap_8
XFILLER_97_431 VDD VSS sg13g2_decap_8
XFILLER_33_0 VDD VSS sg13g2_decap_8
XFILLER_100_904 VDD VSS sg13g2_decap_8
X_2325_ _2325_/RESET_B VSS VDD _2325_/D _2325_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_111_252 VDD VSS sg13g2_decap_8
XFILLER_69_177 VDD VSS sg13g2_decap_8
XFILLER_100_959 VDD VSS sg13g2_decap_8
XFILLER_85_648 VDD VSS sg13g2_fill_1
XFILLER_69_199 VDD VSS sg13g2_fill_1
X_2256_ _2256_/RESET_B VSS VDD _2256_/D _2256_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_38_520 VDD VSS sg13g2_fill_1
X_1207_ VDD _1207_/Y _2251_/Q VSS sg13g2_inv_1
X_2187_ _2187_/RESET_B VSS VDD _2187_/D _2187_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_38_597 VDD VSS sg13g2_decap_8
XFILLER_53_512 VDD VSS sg13g2_decap_4
XFILLER_25_203 VDD VSS sg13g2_decap_8
XFILLER_80_320 VDD VSS sg13g2_decap_8
XFILLER_34_770 VDD VSS sg13g2_decap_8
XFILLER_22_910 VDD VSS sg13g2_decap_8
XFILLER_43_28 VDD VSS sg13g2_decap_8
XFILLER_40_217 VDD VSS sg13g2_decap_8
XFILLER_80_397 VDD VSS sg13g2_decap_8
XFILLER_21_420 VDD VSS sg13g2_decap_8
XFILLER_33_280 VDD VSS sg13g2_decap_8
XFILLER_22_987 VDD VSS sg13g2_decap_8
XFILLER_21_497 VDD VSS sg13g2_decap_8
XFILLER_88_1054 VDD VSS sg13g2_decap_8
XFILLER_111_7 VDD VSS sg13g2_decap_8
XFILLER_107_569 VDD VSS sg13g2_decap_8
XFILLER_108_21 VDD VSS sg13g2_decap_8
XFILLER_49_1049 VDD VSS sg13g2_decap_8
XFILLER_68_14 VDD VSS sg13g2_decap_8
XFILLER_89_943 VDD VSS sg13g2_decap_8
XFILLER_89_965 VDD VSS sg13g2_decap_8
XFILLER_103_742 VDD VSS sg13g2_fill_1
XFILLER_108_98 VDD VSS sg13g2_decap_8
XFILLER_1_847 VDD VSS sg13g2_decap_8
XFILLER_102_241 VDD VSS sg13g2_decap_8
XFILLER_88_464 VDD VSS sg13g2_decap_8
XFILLER_49_818 VDD VSS sg13g2_decap_8
XFILLER_0_357 VDD VSS sg13g2_decap_8
XFILLER_84_35 VDD VSS sg13g2_decap_8
XFILLER_75_147 VDD VSS sg13g2_decap_8
XFILLER_57_873 VDD VSS sg13g2_decap_8
XFILLER_29_553 VDD VSS sg13g2_decap_8
XFILLER_72_821 VDD VSS sg13g2_decap_8
XFILLER_16_203 VDD VSS sg13g2_decap_8
XFILLER_1_1029 VDD VSS sg13g2_decap_8
XFILLER_95_1036 VDD VSS sg13g2_decap_8
X_2178__184 VDD VSS _2178_/RESET_B sg13g2_tiehi
XFILLER_90_139 VDD VSS sg13g2_decap_8
XFILLER_32_707 VDD VSS sg13g2_decap_8
XFILLER_72_898 VDD VSS sg13g2_decap_8
XFILLER_71_364 VDD VSS sg13g2_decap_8
XFILLER_44_578 VDD VSS sg13g2_decap_8
XFILLER_25_770 VDD VSS sg13g2_decap_8
XFILLER_17_84 VDD VSS sg13g2_decap_8
XFILLER_13_910 VDD VSS sg13g2_decap_8
XFILLER_31_217 VDD VSS sg13g2_decap_8
XFILLER_71_397 VDD VSS sg13g2_decap_8
XFILLER_12_420 VDD VSS sg13g2_decap_8
XFILLER_9_903 VDD VSS sg13g2_decap_8
XFILLER_24_280 VDD VSS sg13g2_decap_8
XFILLER_8_413 VDD VSS sg13g2_decap_8
XFILLER_13_987 VDD VSS sg13g2_decap_8
XFILLER_40_795 VDD VSS sg13g2_decap_8
XFILLER_12_497 VDD VSS sg13g2_decap_8
XFILLER_4_630 VDD VSS sg13g2_decap_8
XFILLER_99_729 VDD VSS sg13g2_decap_8
XFILLER_3_140 VDD VSS sg13g2_decap_8
XFILLER_106_580 VDD VSS sg13g2_decap_8
XFILLER_98_239 VDD VSS sg13g2_decap_8
XFILLER_95_924 VDD VSS sg13g2_decap_8
XFILLER_79_475 VDD VSS sg13g2_decap_8
XFILLER_39_317 VDD VSS sg13g2_decap_8
XFILLER_94_412 VDD VSS sg13g2_decap_8
X_2110_ _2110_/A _2110_/B _2110_/Y VDD VSS sg13g2_nor2_1
X_2041_ _2041_/Y _2022_/X _2089_/S _2019_/X _2004_/Y VDD VSS sg13g2_a22oi_1
XFILLER_82_618 VDD VSS sg13g2_decap_8
XFILLER_94_489 VDD VSS sg13g2_decap_8
XFILLER_81_128 VDD VSS sg13g2_decap_8
XFILLER_63_832 VDD VSS sg13g2_decap_8
XFILLER_48_895 VDD VSS sg13g2_fill_1
XFILLER_48_884 VDD VSS sg13g2_fill_1
XFILLER_90_640 VDD VSS sg13g2_decap_8
XFILLER_35_567 VDD VSS sg13g2_decap_8
XFILLER_23_707 VDD VSS sg13g2_decap_8
XFILLER_62_364 VDD VSS sg13g2_fill_2
XFILLER_16_770 VDD VSS sg13g2_decap_8
XFILLER_50_504 VDD VSS sg13g2_decap_8
XFILLER_62_386 VDD VSS sg13g2_decap_8
XFILLER_15_280 VDD VSS sg13g2_decap_8
XFILLER_22_217 VDD VSS sg13g2_decap_8
XFILLER_31_784 VDD VSS sg13g2_decap_8
X_1825_ _1825_/Y _1825_/A _1825_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_294 VDD VSS sg13g2_decap_8
Xhold402 _1334_/Y VDD VSS _1335_/A sg13g2_dlygate4sd3_1
X_1756_ _1761_/B _1756_/B _1763_/A VDD VSS sg13g2_nand2b_1
XFILLER_8_980 VDD VSS sg13g2_decap_8
Xhold435 _2302_/Q VDD VSS hold435/X sg13g2_dlygate4sd3_1
Xhold424 _2305_/Q VDD VSS hold424/X sg13g2_dlygate4sd3_1
Xhold413 _2229_/Q VDD VSS _1416_/A sg13g2_dlygate4sd3_1
XFILLER_7_490 VDD VSS sg13g2_decap_8
Xhold468 _1701_/Y VDD VSS _2315_/D sg13g2_dlygate4sd3_1
XFILLER_104_517 VDD VSS sg13g2_decap_8
X_1687_ _1687_/Y _1724_/S _1693_/A VDD VSS sg13g2_nand2_1
Xhold446 _2207_/Q VDD VSS hold446/X sg13g2_dlygate4sd3_1
Xhold457 _2277_/Q VDD VSS hold457/X sg13g2_dlygate4sd3_1
Xhold479 _2236_/Q VDD VSS hold479/X sg13g2_dlygate4sd3_1
XFILLER_48_1060 VDD VSS sg13g2_fill_1
XFILLER_97_294 VDD VSS sg13g2_decap_8
X_2308_ _2308__81/L_HI VSS VDD _2308_/D _2308_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_58_637 VDD VSS sg13g2_decap_8
XFILLER_38_28 VDD VSS sg13g2_decap_8
XFILLER_86_979 VDD VSS sg13g2_fill_2
XFILLER_57_136 VDD VSS sg13g2_decap_8
XFILLER_94_990 VDD VSS sg13g2_decap_8
XFILLER_85_489 VDD VSS sg13g2_decap_8
X_2239_ _2239_/RESET_B VSS VDD _2239_/D _2239_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_54_843 VDD VSS sg13g2_decap_8
XFILLER_65_191 VDD VSS sg13g2_decap_8
XFILLER_38_383 VDD VSS sg13g2_decap_8
XFILLER_81_673 VDD VSS sg13g2_decap_8
XFILLER_80_150 VDD VSS sg13g2_decap_8
XFILLER_26_567 VDD VSS sg13g2_decap_8
XFILLER_53_375 VDD VSS sg13g2_decap_8
XFILLER_14_707 VDD VSS sg13g2_decap_8
XFILLER_55_1031 VDD VSS sg13g2_decap_8
XFILLER_13_217 VDD VSS sg13g2_decap_8
XFILLER_110_77 VDD VSS sg13g2_decap_8
XFILLER_41_559 VDD VSS sg13g2_fill_1
XFILLER_16_1015 VDD VSS sg13g2_decap_8
XFILLER_22_784 VDD VSS sg13g2_decap_8
XFILLER_10_924 VDD VSS sg13g2_decap_8
XFILLER_103_1029 VDD VSS sg13g2_decap_8
XFILLER_108_801 VDD VSS sg13g2_decap_8
XFILLER_6_917 VDD VSS sg13g2_decap_8
XFILLER_21_294 VDD VSS sg13g2_decap_8
XFILLER_5_427 VDD VSS sg13g2_decap_8
XFILLER_108_878 VDD VSS sg13g2_decap_8
XFILLER_79_35 VDD VSS sg13g2_decap_8
XFILLER_107_388 VDD VSS sg13g2_decap_8
XFILLER_1_644 VDD VSS sg13g2_decap_8
XFILLER_76_401 VDD VSS sg13g2_decap_8
XFILLER_49_615 VDD VSS sg13g2_decap_8
XFILLER_0_154 VDD VSS sg13g2_decap_8
XFILLER_88_283 VDD VSS sg13g2_decap_8
XFILLER_95_56 VDD VSS sg13g2_decap_8
XFILLER_23_1008 VDD VSS sg13g2_decap_8
XFILLER_49_648 VDD VSS sg13g2_decap_8
XFILLER_48_125 VDD VSS sg13g2_decap_8
XFILLER_77_979 VDD VSS sg13g2_decap_8
XFILLER_91_426 VDD VSS sg13g2_decap_8
XFILLER_57_681 VDD VSS sg13g2_decap_8
XFILLER_45_821 VDD VSS sg13g2_decap_8
XFILLER_29_350 VDD VSS sg13g2_decap_8
XFILLER_45_832 VDD VSS sg13g2_fill_1
XFILLER_56_180 VDD VSS sg13g2_decap_8
XFILLER_72_662 VDD VSS sg13g2_fill_1
XFILLER_60_813 VDD VSS sg13g2_decap_8
XFILLER_45_876 VDD VSS sg13g2_fill_1
XFILLER_17_567 VDD VSS sg13g2_decap_8
XFILLER_32_504 VDD VSS sg13g2_decap_8
XFILLER_44_364 VDD VSS sg13g2_decap_8
XFILLER_71_183 VDD VSS sg13g2_decap_8
XFILLER_60_879 VDD VSS sg13g2_decap_8
XFILLER_9_700 VDD VSS sg13g2_decap_8
XFILLER_8_210 VDD VSS sg13g2_decap_8
XFILLER_13_784 VDD VSS sg13g2_decap_8
XFILLER_74_7 VDD VSS sg13g2_decap_8
XFILLER_40_592 VDD VSS sg13g2_decap_8
XFILLER_12_294 VDD VSS sg13g2_decap_8
XFILLER_9_777 VDD VSS sg13g2_decap_8
XFILLER_8_287 VDD VSS sg13g2_decap_8
X_1610_ _1639_/A _1610_/B _1610_/Y VDD VSS sg13g2_nor2_1
XFILLER_5_21 VDD VSS sg13g2_decap_8
XFILLER_99_504 VDD VSS sg13g2_decap_4
X_1541_ _1576_/A _1541_/B _2276_/D VDD VSS sg13g2_nor2_1
XFILLER_5_994 VDD VSS sg13g2_decap_8
XFILLER_99_548 VDD VSS sg13g2_decap_8
X_1472_ _1602_/B VDD _1472_/Y VSS _1376_/A _1479_/A2 sg13g2_o21ai_1
XFILLER_5_98 VDD VSS sg13g2_decap_8
XFILLER_86_209 VDD VSS sg13g2_decap_8
XFILLER_79_250 VDD VSS sg13g2_decap_8
XFILLER_67_401 VDD VSS sg13g2_decap_8
XFILLER_95_721 VDD VSS sg13g2_fill_2
XFILLER_55_607 VDD VSS sg13g2_fill_1
XFILLER_39_147 VDD VSS sg13g2_decap_8
XFILLER_95_787 VDD VSS sg13g2_decap_8
XFILLER_82_415 VDD VSS sg13g2_decap_8
XFILLER_67_478 VDD VSS sg13g2_decap_8
XFILLER_54_106 VDD VSS sg13g2_decap_8
XFILLER_78_1042 VDD VSS sg13g2_decap_8
X_2024_ _2022_/S _1999_/A _1901_/B _1931_/A _1914_/A _2021_/S _2024_/X VDD VSS sg13g2_mux4_1
XFILLER_36_854 VDD VSS sg13g2_decap_8
XFILLER_47_191 VDD VSS sg13g2_decap_8
XFILLER_39_1004 VDD VSS sg13g2_decap_8
XFILLER_23_504 VDD VSS sg13g2_decap_8
XFILLER_35_364 VDD VSS sg13g2_decap_8
XFILLER_63_684 VDD VSS sg13g2_decap_4
XFILLER_51_835 VDD VSS sg13g2_decap_4
XFILLER_50_367 VDD VSS sg13g2_decap_8
XFILLER_31_581 VDD VSS sg13g2_decap_8
XFILLER_109_609 VDD VSS sg13g2_decap_8
X_1808_ _1797_/Y VDD _1825_/B VSS _1823_/A _1823_/B sg13g2_o21ai_1
XFILLER_108_119 VDD VSS sg13g2_decap_8
XFILLER_105_826 VDD VSS sg13g2_decap_8
XFILLER_104_314 VDD VSS sg13g2_decap_8
X_1739_ VDD VSS _1767_/B _1728_/Y _1898_/A _1727_/Y _1763_/A _1729_/Y sg13g2_a221oi_1
XFILLER_85_1057 VDD VSS sg13g2_decap_4
XFILLER_49_49 VDD VSS sg13g2_decap_8
Xhold298 _1226_/X VDD VSS _2358_/D sg13g2_dlygate4sd3_1
XFILLER_98_581 VDD VSS sg13g2_decap_8
XFILLER_59_957 VDD VSS sg13g2_decap_8
XFILLER_100_553 VDD VSS sg13g2_fill_2
XFILLER_74_905 VDD VSS sg13g2_decap_8
XFILLER_100_531 VDD VSS sg13g2_decap_8
XFILLER_85_231 VDD VSS sg13g2_decap_8
XFILLER_46_607 VDD VSS sg13g2_decap_8
XFILLER_105_77 VDD VSS sg13g2_decap_8
XFILLER_27_854 VDD VSS sg13g2_decap_8
XFILLER_45_139 VDD VSS sg13g2_decap_8
XFILLER_14_504 VDD VSS sg13g2_decap_8
XFILLER_53_150 VDD VSS sg13g2_fill_1
XFILLER_26_364 VDD VSS sg13g2_decap_8
XFILLER_81_14 VDD VSS sg13g2_decap_8
XFILLER_41_301 VDD VSS sg13g2_decap_8
XFILLER_42_868 VDD VSS sg13g2_decap_8
XFILLER_14_63 VDD VSS sg13g2_decap_8
XFILLER_22_581 VDD VSS sg13g2_decap_8
XFILLER_10_721 VDD VSS sg13g2_decap_8
XFILLER_6_714 VDD VSS sg13g2_decap_8
XFILLER_5_224 VDD VSS sg13g2_decap_8
XFILLER_10_798 VDD VSS sg13g2_decap_8
XFILLER_108_675 VDD VSS sg13g2_decap_8
XFILLER_100_0 VDD VSS sg13g2_decap_8
XFILLER_2_931 VDD VSS sg13g2_decap_8
XFILLER_30_84 VDD VSS sg13g2_decap_8
XFILLER_96_507 VDD VSS sg13g2_decap_8
XFILLER_1_441 VDD VSS sg13g2_decap_8
XFILLER_49_412 VDD VSS sg13g2_decap_8
XFILLER_65_916 VDD VSS sg13g2_decap_8
XFILLER_7_1057 VDD VSS sg13g2_decap_4
XFILLER_92_735 VDD VSS sg13g2_decap_8
XFILLER_76_275 VDD VSS sg13g2_decap_8
XFILLER_49_489 VDD VSS sg13g2_fill_2
XFILLER_49_478 VDD VSS sg13g2_decap_8
XFILLER_80_908 VDD VSS sg13g2_decap_4
XFILLER_91_234 VDD VSS sg13g2_decap_8
XFILLER_18_854 VDD VSS sg13g2_decap_8
XFILLER_45_651 VDD VSS sg13g2_fill_1
XFILLER_17_364 VDD VSS sg13g2_decap_8
XFILLER_55_70 VDD VSS sg13g2_fill_2
XFILLER_32_301 VDD VSS sg13g2_decap_8
XFILLER_60_654 VDD VSS sg13g2_fill_1
XFILLER_33_868 VDD VSS sg13g2_decap_8
XFILLER_20_518 VDD VSS sg13g2_decap_8
XFILLER_32_378 VDD VSS sg13g2_decap_8
XFILLER_71_80 VDD VSS sg13g2_decap_4
XFILLER_13_581 VDD VSS sg13g2_decap_8
XFILLER_9_574 VDD VSS sg13g2_decap_8
XFILLER_5_791 VDD VSS sg13g2_decap_8
X_1524_ _1524_/Y _1589_/C _1584_/B VDD VSS sg13g2_nand2_1
XFILLER_102_818 VDD VSS sg13g2_decap_8
XFILLER_99_367 VDD VSS sg13g2_fill_1
XFILLER_87_507 VDD VSS sg13g2_decap_8
X_1455_ _1455_/A _1455_/B _1455_/Y VDD VSS sg13g2_nor2_1
XFILLER_45_1052 VDD VSS sg13g2_decap_8
XFILLER_110_851 VDD VSS sg13g2_decap_8
X_1386_ _1386_/Y _1386_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_55_459 VDD VSS sg13g2_decap_8
X_2007_ _2071_/A _2007_/B _2037_/A VDD VSS sg13g2_and2_1
XFILLER_82_278 VDD VSS sg13g2_decap_8
XFILLER_70_407 VDD VSS sg13g2_decap_8
XFILLER_36_651 VDD VSS sg13g2_decap_8
XFILLER_64_993 VDD VSS sg13g2_decap_8
XFILLER_35_161 VDD VSS sg13g2_decap_8
XFILLER_23_301 VDD VSS sg13g2_decap_8
XFILLER_51_654 VDD VSS sg13g2_decap_8
XFILLER_24_868 VDD VSS sg13g2_decap_8
XFILLER_50_120 VDD VSS sg13g2_decap_8
XFILLER_11_518 VDD VSS sg13g2_decap_8
XFILLER_23_378 VDD VSS sg13g2_decap_8
XFILLER_109_406 VDD VSS sg13g2_decap_8
XFILLER_52_1045 VDD VSS sg13g2_decap_8
XFILLER_13_1029 VDD VSS sg13g2_decap_8
XFILLER_3_728 VDD VSS sg13g2_decap_8
XFILLER_105_623 VDD VSS sg13g2_decap_8
XFILLER_2_238 VDD VSS sg13g2_decap_8
XFILLER_4_7 VDD VSS sg13g2_decap_8
XFILLER_104_133 VDD VSS sg13g2_decap_8
XFILLER_104_188 VDD VSS sg13g2_decap_8
XFILLER_78_529 VDD VSS sg13g2_decap_8
XFILLER_76_14 VDD VSS sg13g2_decap_8
XFILLER_59_721 VDD VSS sg13g2_decap_8
XFILLER_101_851 VDD VSS sg13g2_decap_8
XFILLER_86_584 VDD VSS sg13g2_decap_8
XFILLER_74_702 VDD VSS sg13g2_decap_8
XFILLER_73_201 VDD VSS sg13g2_decap_8
XFILLER_92_35 VDD VSS sg13g2_decap_8
XFILLER_27_651 VDD VSS sg13g2_decap_8
XFILLER_61_418 VDD VSS sg13g2_decap_8
XFILLER_54_481 VDD VSS sg13g2_decap_8
XFILLER_14_301 VDD VSS sg13g2_decap_8
XFILLER_26_161 VDD VSS sg13g2_decap_8
XFILLER_70_941 VDD VSS sg13g2_decap_8
XFILLER_42_665 VDD VSS sg13g2_decap_8
XFILLER_30_805 VDD VSS sg13g2_decap_8
XFILLER_15_868 VDD VSS sg13g2_decap_8
XFILLER_109_1057 VDD VSS sg13g2_decap_4
XFILLER_14_378 VDD VSS sg13g2_decap_8
XFILLER_25_84 VDD VSS sg13g2_decap_8
XFILLER_6_511 VDD VSS sg13g2_decap_8
XFILLER_10_595 VDD VSS sg13g2_decap_8
XFILLER_109_973 VDD VSS sg13g2_decap_8
XFILLER_108_450 VDD VSS sg13g2_decap_8
XFILLER_6_588 VDD VSS sg13g2_decap_8
XFILLER_29_1036 VDD VSS sg13g2_decap_8
XFILLER_111_637 VDD VSS sg13g2_decap_8
X_2340__143 VDD VSS _2340_/RESET_B sg13g2_tiehi
XFILLER_96_315 VDD VSS sg13g2_decap_8
XFILLER_37_7 VDD VSS sg13g2_decap_8
XFILLER_77_551 VDD VSS sg13g2_decap_8
XFILLER_110_147 VDD VSS sg13g2_decap_8
XFILLER_38_905 VDD VSS sg13g2_decap_8
X_1240_ _1248_/B _2295_/Q _2257_/Q VDD VSS sg13g2_xnor2_1
XFILLER_65_724 VDD VSS sg13g2_decap_8
XFILLER_2_77 VDD VSS sg13g2_decap_8
XFILLER_49_253 VDD VSS sg13g2_decap_8
XFILLER_64_212 VDD VSS sg13g2_decap_8
XFILLER_37_448 VDD VSS sg13g2_decap_8
XFILLER_92_565 VDD VSS sg13g2_decap_8
XFILLER_18_651 VDD VSS sg13g2_decap_8
XFILLER_66_91 VDD VSS sg13g2_decap_8
XFILLER_75_1023 VDD VSS sg13g2_fill_2
XFILLER_46_982 VDD VSS sg13g2_decap_8
XFILLER_17_161 VDD VSS sg13g2_decap_8
XFILLER_33_665 VDD VSS sg13g2_decap_8
XFILLER_21_805 VDD VSS sg13g2_decap_8
XFILLER_36_1029 VDD VSS sg13g2_decap_8
XFILLER_20_315 VDD VSS sg13g2_decap_8
XFILLER_60_484 VDD VSS sg13g2_decap_4
XFILLER_32_175 VDD VSS sg13g2_decap_8
XFILLER_9_371 VDD VSS sg13g2_decap_8
XFILLER_63_0 VDD VSS sg13g2_decap_8
XFILLER_82_1005 VDD VSS sg13g2_decap_8
XFILLER_88_816 VDD VSS sg13g2_decap_8
XFILLER_102_637 VDD VSS sg13g2_fill_2
X_1507_ _1507_/A _1514_/A _1507_/Y VDD VSS sg13g2_nor2_1
X_1438_ _1439_/A _1429_/Y hold452/X _1429_/B _1379_/A VDD VSS sg13g2_a22oi_1
XFILLER_87_337 VDD VSS sg13g2_decap_8
XFILLER_101_147 VDD VSS sg13g2_decap_4
XFILLER_96_871 VDD VSS sg13g2_decap_8
XFILLER_29_938 VDD VSS sg13g2_decap_8
XFILLER_68_551 VDD VSS sg13g2_decap_8
XFILLER_83_543 VDD VSS sg13g2_decap_8
XFILLER_95_392 VDD VSS sg13g2_decap_8
X_1369_ _1368_/Y VDD _2211_/D VSS _1364_/Y _1367_/B sg13g2_o21ai_1
XFILLER_56_735 VDD VSS sg13g2_decap_8
XFILLER_46_28 VDD VSS sg13g2_decap_8
XFILLER_28_448 VDD VSS sg13g2_decap_8
XFILLER_55_245 VDD VSS sg13g2_decap_8
XFILLER_71_727 VDD VSS sg13g2_decap_8
XFILLER_70_248 VDD VSS sg13g2_decap_8
XFILLER_102_56 VDD VSS sg13g2_decap_8
XFILLER_24_665 VDD VSS sg13g2_decap_8
XFILLER_12_805 VDD VSS sg13g2_decap_8
XFILLER_62_49 VDD VSS sg13g2_decap_8
XFILLER_11_315 VDD VSS sg13g2_decap_8
XFILLER_23_175 VDD VSS sg13g2_decap_8
XFILLER_109_203 VDD VSS sg13g2_decap_8
XFILLER_7_308 VDD VSS sg13g2_decap_8
XFILLER_109_247 VDD VSS sg13g2_decap_8
XFILLER_20_882 VDD VSS sg13g2_decap_8
XIO_BOND_in_ready_pad in_ready_PAD bondpad_70x70
XFILLER_11_42 VDD VSS sg13g2_decap_8
XFILLER_3_525 VDD VSS sg13g2_decap_8
XFILLER_106_965 VDD VSS sg13g2_decap_8
XFILLER_105_442 VDD VSS sg13g2_decap_8
XFILLER_105_497 VDD VSS sg13g2_fill_2
XFILLER_87_35 VDD VSS sg13g2_decap_8
XFILLER_87_871 VDD VSS sg13g2_decap_8
XFILLER_98_1012 VDD VSS sg13g2_fill_2
XFILLER_101_692 VDD VSS sg13g2_decap_8
XFILLER_86_370 VDD VSS sg13g2_decap_8
XFILLER_47_757 VDD VSS sg13g2_decap_8
XFILLER_19_448 VDD VSS sg13g2_decap_8
XFILLER_100_191 VDD VSS sg13g2_decap_8
XFILLER_46_245 VDD VSS sg13g2_decap_8
XFILLER_46_234 VDD VSS sg13g2_decap_8
XFILLER_55_790 VDD VSS sg13g2_decap_8
XFILLER_61_259 VDD VSS sg13g2_decap_8
XFILLER_42_440 VDD VSS sg13g2_decap_8
XFILLER_43_996 VDD VSS sg13g2_decap_8
XFILLER_30_602 VDD VSS sg13g2_decap_8
XFILLER_15_665 VDD VSS sg13g2_decap_8
XFILLER_14_175 VDD VSS sg13g2_decap_8
XFILLER_30_679 VDD VSS sg13g2_decap_8
XFILLER_52_82 VDD VSS sg13g2_decap_8
XFILLER_11_882 VDD VSS sg13g2_decap_8
XFILLER_109_770 VDD VSS sg13g2_decap_8
X_2188__164 VDD VSS _2188_/RESET_B sg13g2_tiehi
XFILLER_10_392 VDD VSS sg13g2_decap_8
XFILLER_7_875 VDD VSS sg13g2_decap_8
XFILLER_6_385 VDD VSS sg13g2_decap_8
XFILLER_108_291 VDD VSS sg13g2_decap_8
XFILLER_112_924 VDD VSS sg13g2_decap_8
X_2341_ _2341_/RESET_B VSS VDD _2341_/D _2341_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_96_112 VDD VSS sg13g2_decap_8
XFILLER_97_668 VDD VSS sg13g2_decap_8
XFILLER_111_434 VDD VSS sg13g2_decap_8
XFILLER_69_348 VDD VSS sg13g2_decap_8
X_2299__115 VDD VSS _2299_/RESET_B sg13g2_tiehi
X_2272_ _2272_/RESET_B VSS VDD _2272_/D _2272_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_42_1022 VDD VSS sg13g2_decap_8
X_1223_ _2150_/A _2150_/B _2362_/D VDD VSS sg13g2_and2_1
XFILLER_38_702 VDD VSS sg13g2_decap_8
XFILLER_96_189 VDD VSS sg13g2_decap_8
XFILLER_93_852 VDD VSS sg13g2_decap_8
XFILLER_92_340 VDD VSS sg13g2_decap_8
XFILLER_65_543 VDD VSS sg13g2_decap_8
XFILLER_38_779 VDD VSS sg13g2_decap_8
XFILLER_37_245 VDD VSS sg13g2_decap_8
XFILLER_80_502 VDD VSS sg13g2_decap_8
XFILLER_65_598 VDD VSS sg13g2_decap_8
XFILLER_53_738 VDD VSS sg13g2_decap_4
XFILLER_52_226 VDD VSS sg13g2_fill_1
XFILLER_34_952 VDD VSS sg13g2_decap_8
XFILLER_21_602 VDD VSS sg13g2_decap_8
XFILLER_33_462 VDD VSS sg13g2_decap_8
XFILLER_60_270 VDD VSS sg13g2_decap_8
XFILLER_20_112 VDD VSS sg13g2_decap_8
X_1987_ _1988_/B _1987_/A _1987_/B VDD VSS sg13g2_xnor2_1
XFILLER_21_679 VDD VSS sg13g2_decap_8
XFILLER_20_189 VDD VSS sg13g2_decap_8
XFILLER_106_217 VDD VSS sg13g2_decap_8
XFILLER_103_924 VDD VSS sg13g2_decap_8
XFILLER_88_635 VDD VSS sg13g2_decap_8
XFILLER_87_123 VDD VSS sg13g2_fill_2
XFILLER_0_539 VDD VSS sg13g2_decap_8
XFILLER_88_679 VDD VSS sg13g2_decap_8
XFILLER_102_456 VDD VSS sg13g2_decap_8
XFILLER_57_38 VDD VSS sg13g2_fill_1
XFILLER_29_735 VDD VSS sg13g2_decap_8
XFILLER_28_245 VDD VSS sg13g2_decap_8
XFILLER_84_885 VDD VSS sg13g2_decap_8
XFILLER_71_502 VDD VSS sg13g2_decap_8
XFILLER_71_557 VDD VSS sg13g2_decap_8
X_2254__243 VDD VSS _2254_/RESET_B sg13g2_tiehi
XFILLER_25_952 VDD VSS sg13g2_decap_8
XFILLER_43_237 VDD VSS sg13g2_decap_8
XFILLER_40_900 VDD VSS sg13g2_decap_8
XFILLER_12_602 VDD VSS sg13g2_decap_8
XFILLER_24_462 VDD VSS sg13g2_decap_8
XFILLER_11_112 VDD VSS sg13g2_decap_8
XFILLER_19_1057 VDD VSS sg13g2_decap_4
XFILLER_106_1049 VDD VSS sg13g2_decap_8
XFILLER_40_977 VDD VSS sg13g2_decap_8
XFILLER_7_105 VDD VSS sg13g2_decap_8
XFILLER_12_679 VDD VSS sg13g2_decap_8
XFILLER_11_189 VDD VSS sg13g2_decap_8
XFILLER_22_63 VDD VSS sg13g2_decap_8
XFILLER_4_812 VDD VSS sg13g2_decap_8
XFILLER_98_56 VDD VSS sg13g2_decap_8
XFILLER_3_322 VDD VSS sg13g2_decap_8
XFILLER_106_762 VDD VSS sg13g2_decap_8
XFILLER_79_624 VDD VSS sg13g2_decap_8
XFILLER_65_1022 VDD VSS sg13g2_decap_8
XFILLER_4_889 VDD VSS sg13g2_decap_8
XFILLER_79_657 VDD VSS sg13g2_decap_8
XFILLER_78_112 VDD VSS sg13g2_decap_8
XFILLER_3_399 VDD VSS sg13g2_decap_8
XFILLER_75_841 VDD VSS sg13g2_decap_8
XFILLER_66_329 VDD VSS sg13g2_decap_8
XFILLER_19_245 VDD VSS sg13g2_decap_8
XFILLER_74_373 VDD VSS sg13g2_fill_1
XFILLER_47_576 VDD VSS sg13g2_decap_8
XFILLER_47_587 VDD VSS sg13g2_fill_2
XFILLER_35_749 VDD VSS sg13g2_decap_8
XFILLER_16_952 VDD VSS sg13g2_decap_8
XFILLER_72_1004 VDD VSS sg13g2_decap_8
XFILLER_90_888 VDD VSS sg13g2_decap_8
XFILLER_62_568 VDD VSS sg13g2_fill_2
XFILLER_15_462 VDD VSS sg13g2_decap_8
XFILLER_34_259 VDD VSS sg13g2_decap_8
X_1910_ _1943_/B _1943_/A _1911_/B VDD VSS sg13g2_nor2b_1
XFILLER_43_793 VDD VSS sg13g2_decap_8
X_1841_ _1934_/B _2245_/Q _2204_/Q VDD VSS sg13g2_xnor2_1
XFILLER_31_966 VDD VSS sg13g2_decap_8
XFILLER_8_21 VDD VSS sg13g2_decap_8
XFILLER_30_476 VDD VSS sg13g2_decap_8
X_1772_ _1877_/B _1772_/A _1772_/B VDD VSS sg13g2_xnor2_1
XFILLER_8_98 VDD VSS sg13g2_decap_8
Xin_data_pads\[5\].in_data_pad IOVDD IOVSS _1382_/A in_data_PADs[5] VDD VSS sg13g2_IOPadIn
XFILLER_7_672 VDD VSS sg13g2_decap_8
XFILLER_6_182 VDD VSS sg13g2_decap_8
XFILLER_112_721 VDD VSS sg13g2_decap_8
X_2324_ _2324_/RESET_B VSS VDD _2324_/D _2324_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_97_421 VDD VSS sg13g2_fill_2
XFILLER_69_134 VDD VSS sg13g2_decap_8
XFILLER_98_999 VDD VSS sg13g2_fill_1
XFILLER_111_231 VDD VSS sg13g2_decap_8
XFILLER_69_156 VDD VSS sg13g2_decap_8
XFILLER_26_0 VDD VSS sg13g2_decap_8
XFILLER_112_798 VDD VSS sg13g2_decap_8
XFILLER_78_690 VDD VSS sg13g2_decap_8
XFILLER_84_126 VDD VSS sg13g2_fill_2
X_2255_ _2255_/RESET_B VSS VDD _2255_/D _2255_/Q clkload4/A sg13g2_dfrbpq_1
X_1206_ VDD _1206_/Y _2271_/Q VSS sg13g2_inv_1
X_2186_ _2186_/RESET_B VSS VDD _2186_/D _2186_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_38_576 VDD VSS sg13g2_decap_8
XFILLER_92_192 VDD VSS sg13g2_decap_8
XFILLER_26_749 VDD VSS sg13g2_decap_8
XFILLER_53_535 VDD VSS sg13g2_fill_1
XFILLER_80_376 VDD VSS sg13g2_decap_8
XFILLER_25_259 VDD VSS sg13g2_decap_8
XFILLER_61_590 VDD VSS sg13g2_decap_8
XFILLER_22_966 VDD VSS sg13g2_decap_8
XFILLER_21_476 VDD VSS sg13g2_decap_8
XFILLER_88_1000 VDD VSS sg13g2_decap_8
XFILLER_5_609 VDD VSS sg13g2_decap_8
XFILLER_49_1006 VDD VSS sg13g2_fill_2
XFILLER_4_119 VDD VSS sg13g2_decap_8
XFILLER_107_548 VDD VSS sg13g2_decap_8
XFILLER_104_7 VDD VSS sg13g2_decap_8
XFILLER_89_922 VDD VSS sg13g2_decap_8
XFILLER_108_77 VDD VSS sg13g2_decap_8
XFILLER_1_826 VDD VSS sg13g2_decap_8
XFILLER_88_443 VDD VSS sg13g2_decap_8
XFILLER_0_336 VDD VSS sg13g2_decap_8
XFILLER_103_798 VDD VSS sg13g2_decap_4
XFILLER_75_126 VDD VSS sg13g2_decap_8
XFILLER_25_1050 VDD VSS sg13g2_decap_8
XFILLER_48_329 VDD VSS sg13g2_decap_8
XFILLER_84_14 VDD VSS sg13g2_decap_8
XFILLER_56_340 VDD VSS sg13g2_decap_8
XFILLER_29_532 VDD VSS sg13g2_decap_8
XFILLER_95_1015 VDD VSS sg13g2_decap_8
XFILLER_90_129 VDD VSS sg13g2_decap_4
XFILLER_1_1008 VDD VSS sg13g2_decap_8
XFILLER_83_192 VDD VSS sg13g2_decap_8
XFILLER_44_557 VDD VSS sg13g2_decap_8
XFILLER_56_384 VDD VSS sg13g2_decap_8
XFILLER_17_63 VDD VSS sg13g2_decap_8
XFILLER_17_749 VDD VSS sg13g2_decap_8
XFILLER_16_259 VDD VSS sg13g2_decap_8
XFILLER_52_590 VDD VSS sg13g2_decap_4
XFILLER_13_966 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[1\].out_data_pad out_data_PADs[1] bondpad_70x70
XFILLER_40_774 VDD VSS sg13g2_decap_8
XFILLER_12_476 VDD VSS sg13g2_decap_8
XFILLER_9_959 VDD VSS sg13g2_decap_8
XFILLER_33_84 VDD VSS sg13g2_decap_8
XFILLER_32_1043 VDD VSS sg13g2_decap_8
XFILLER_8_469 VDD VSS sg13g2_decap_8
XFILLER_99_708 VDD VSS sg13g2_decap_8
XFILLER_98_218 VDD VSS sg13g2_decap_8
XFILLER_4_686 VDD VSS sg13g2_decap_8
XFILLER_3_196 VDD VSS sg13g2_decap_8
XFILLER_95_903 VDD VSS sg13g2_decap_8
XFILLER_79_454 VDD VSS sg13g2_decap_8
XFILLER_67_649 VDD VSS sg13g2_fill_2
XFILLER_66_126 VDD VSS sg13g2_decap_8
X_2040_ _2040_/Y _2040_/A _2149_/A VDD VSS sg13g2_nand2_1
XFILLER_94_468 VDD VSS sg13g2_decap_8
XFILLER_48_863 VDD VSS sg13g2_decap_8
XFILLER_63_811 VDD VSS sg13g2_decap_8
XFILLER_75_693 VDD VSS sg13g2_decap_8
XFILLER_35_546 VDD VSS sg13g2_decap_8
XFILLER_74_91 VDD VSS sg13g2_decap_8
XFILLER_63_888 VDD VSS sg13g2_decap_8
XFILLER_90_696 VDD VSS sg13g2_decap_8
XFILLER_43_590 VDD VSS sg13g2_decap_8
XFILLER_31_763 VDD VSS sg13g2_decap_8
XFILLER_30_273 VDD VSS sg13g2_decap_8
X_1824_ _1930_/A VDD _1826_/A VSS _1822_/B _1878_/B sg13g2_o21ai_1
XIO_FILL_IO_SOUTH_0_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
X_1755_ _1754_/Y VDD _1760_/B VSS _1763_/A _1750_/Y sg13g2_o21ai_1
Xhold436 _1657_/Y VDD VSS _1658_/B sg13g2_dlygate4sd3_1
Xhold425 _1666_/Y VDD VSS _1667_/B sg13g2_dlygate4sd3_1
Xhold414 _2231_/Q VDD VSS _1420_/A sg13g2_dlygate4sd3_1
Xhold403 _2360_/Q VDD VSS _2150_/B sg13g2_dlygate4sd3_1
XFILLER_89_207 VDD VSS sg13g2_decap_8
Xhold447 _2237_/Q VDD VSS hold447/X sg13g2_dlygate4sd3_1
Xhold469 _2235_/Q VDD VSS hold469/X sg13g2_dlygate4sd3_1
X_1686_ _1693_/A _1723_/A _1686_/B VDD VSS sg13g2_xnor2_1
Xhold458 _1547_/Y VDD VSS _1548_/B sg13g2_dlygate4sd3_1
XFILLER_98_785 VDD VSS sg13g2_decap_8
XFILLER_58_616 VDD VSS sg13g2_decap_8
XFILLER_86_958 VDD VSS sg13g2_decap_8
XFILLER_112_595 VDD VSS sg13g2_decap_8
XFILLER_100_724 VDD VSS sg13g2_decap_8
XFILLER_97_284 VDD VSS sg13g2_decap_4
X_2307_ _2307__83/L_HI VSS VDD _2307_/D _2307_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_57_115 VDD VSS sg13g2_decap_8
XFILLER_100_779 VDD VSS sg13g2_decap_8
X_2238_ _2238_/RESET_B VSS VDD _2238_/D _2238_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_54_822 VDD VSS sg13g2_decap_8
XFILLER_39_885 VDD VSS sg13g2_decap_8
XFILLER_38_362 VDD VSS sg13g2_decap_8
X_2169_ _2169_/RESET_B VSS VDD _2169_/D _2169_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_93_490 VDD VSS sg13g2_fill_2
XFILLER_66_693 VDD VSS sg13g2_decap_8
XFILLER_26_546 VDD VSS sg13g2_decap_8
XFILLER_65_170 VDD VSS sg13g2_decap_8
XFILLER_53_310 VDD VSS sg13g2_fill_2
XFILLER_54_28 VDD VSS sg13g2_decap_8
XFILLER_81_652 VDD VSS sg13g2_decap_8
XFILLER_54_899 VDD VSS sg13g2_decap_8
XFILLER_41_516 VDD VSS sg13g2_decap_8
XFILLER_110_56 VDD VSS sg13g2_decap_8
XFILLER_22_763 VDD VSS sg13g2_decap_8
XFILLER_10_903 VDD VSS sg13g2_decap_8
XFILLER_103_1008 VDD VSS sg13g2_decap_8
XFILLER_70_49 VDD VSS sg13g2_decap_8
XFILLER_21_273 VDD VSS sg13g2_decap_8
XFILLER_107_312 VDD VSS sg13g2_decap_8
XFILLER_5_406 VDD VSS sg13g2_decap_8
XFILLER_108_857 VDD VSS sg13g2_decap_8
XFILLER_107_323 VDD VSS sg13g2_fill_1
XFILLER_79_14 VDD VSS sg13g2_decap_8
XFILLER_1_623 VDD VSS sg13g2_decap_8
XFILLER_103_551 VDD VSS sg13g2_decap_4
XFILLER_0_133 VDD VSS sg13g2_decap_8
XFILLER_77_958 VDD VSS sg13g2_decap_8
XFILLER_103_595 VDD VSS sg13g2_decap_8
XFILLER_88_262 VDD VSS sg13g2_decap_8
XFILLER_95_35 VDD VSS sg13g2_decap_8
XFILLER_49_638 VDD VSS sg13g2_fill_1
XFILLER_48_104 VDD VSS sg13g2_decap_8
XFILLER_92_906 VDD VSS sg13g2_fill_2
XFILLER_92_939 VDD VSS sg13g2_decap_8
XFILLER_85_980 VDD VSS sg13g2_decap_8
XFILLER_85_991 VDD VSS sg13g2_fill_2
XFILLER_57_660 VDD VSS sg13g2_decap_8
XFILLER_28_84 VDD VSS sg13g2_decap_8
XFILLER_63_118 VDD VSS sg13g2_decap_8
XFILLER_72_641 VDD VSS sg13g2_decap_8
XFILLER_17_546 VDD VSS sg13g2_decap_8
XFILLER_44_343 VDD VSS sg13g2_decap_8
XFILLER_71_162 VDD VSS sg13g2_decap_8
XFILLER_60_858 VDD VSS sg13g2_decap_8
XFILLER_40_571 VDD VSS sg13g2_decap_8
XFILLER_13_763 VDD VSS sg13g2_decap_8
XFILLER_12_273 VDD VSS sg13g2_decap_8
XFILLER_9_756 VDD VSS sg13g2_decap_8
XFILLER_8_266 VDD VSS sg13g2_decap_8
XFILLER_67_7 VDD VSS sg13g2_decap_8
X_1540_ _1540_/Y _1527_/Y _1539_/Y hold475/X _1527_/B VDD VSS sg13g2_a22oi_1
XFILLER_99_527 VDD VSS sg13g2_decap_8
XFILLER_5_973 VDD VSS sg13g2_decap_8
X_1471_ VSS VDD _1199_/Y _1479_/A2 _2254_/D _1470_/Y sg13g2_a21oi_1
XFILLER_4_483 VDD VSS sg13g2_decap_8
XFILLER_5_77 VDD VSS sg13g2_decap_8
XFILLER_95_700 VDD VSS sg13g2_decap_8
XFILLER_94_210 VDD VSS sg13g2_decap_8
XFILLER_79_284 VDD VSS sg13g2_fill_2
XFILLER_95_766 VDD VSS sg13g2_decap_8
XFILLER_83_906 VDD VSS sg13g2_decap_8
XFILLER_67_457 VDD VSS sg13g2_decap_8
XFILLER_39_126 VDD VSS sg13g2_decap_8
XFILLER_94_254 VDD VSS sg13g2_decap_8
XFILLER_78_1021 VDD VSS sg13g2_decap_8
XFILLER_76_991 VDD VSS sg13g2_decap_8
X_2023_ _2022_/X _2074_/A _2020_/Y _2323_/D VDD VSS sg13g2_a21o_1
XFILLER_36_833 VDD VSS sg13g2_decap_8
XFILLER_91_983 VDD VSS sg13g2_fill_2
XFILLER_63_663 VDD VSS sg13g2_decap_8
XFILLER_51_814 VDD VSS sg13g2_decap_8
XFILLER_35_343 VDD VSS sg13g2_decap_8
X_2350__101 VDD VSS _2350_/RESET_B sg13g2_tiehi
XFILLER_62_162 VDD VSS sg13g2_decap_8
X_2170__200 VDD VSS _2170_/RESET_B sg13g2_tiehi
XFILLER_93_0 VDD VSS sg13g2_decap_8
XFILLER_50_346 VDD VSS sg13g2_fill_2
XFILLER_31_560 VDD VSS sg13g2_decap_8
X_1807_ _1795_/A VDD _1823_/B VSS _1801_/Y _1806_/Y sg13g2_o21ai_1
XFILLER_102_1041 VDD VSS sg13g2_decap_8
XFILLER_85_1003 VDD VSS sg13g2_fill_1
XFILLER_85_1036 VDD VSS sg13g2_decap_8
XFILLER_105_805 VDD VSS sg13g2_decap_8
X_1738_ _1898_/B _1915_/B _1767_/B VDD VSS sg13g2_and2_1
X_1669_ _1669_/Y _1646_/Y _1668_/X hold422/X _1189_/Y VDD VSS sg13g2_a22oi_1
XFILLER_49_28 VDD VSS sg13g2_decap_8
XFILLER_98_560 VDD VSS sg13g2_decap_8
XFILLER_86_700 VDD VSS sg13g2_decap_8
Xhold299 _2354_/Q VDD VSS _1220_/A sg13g2_dlygate4sd3_1
XFILLER_86_711 VDD VSS sg13g2_fill_1
XFILLER_100_510 VDD VSS sg13g2_decap_8
XFILLER_85_210 VDD VSS sg13g2_decap_8
XFILLER_59_936 VDD VSS sg13g2_decap_8
XFILLER_58_413 VDD VSS sg13g2_fill_2
XFILLER_112_392 VDD VSS sg13g2_decap_8
XFILLER_105_56 VDD VSS sg13g2_decap_8
XFILLER_86_788 VDD VSS sg13g2_decap_8
XFILLER_65_49 VDD VSS sg13g2_decap_8
XFILLER_39_682 VDD VSS sg13g2_decap_8
XFILLER_27_833 VDD VSS sg13g2_decap_8
XFILLER_26_343 VDD VSS sg13g2_decap_8
XFILLER_81_482 VDD VSS sg13g2_decap_8
XFILLER_42_847 VDD VSS sg13g2_decap_8
XFILLER_50_880 VDD VSS sg13g2_decap_8
XFILLER_22_560 VDD VSS sg13g2_decap_8
XFILLER_14_42 VDD VSS sg13g2_decap_8
XFILLER_10_700 VDD VSS sg13g2_decap_8
XFILLER_5_203 VDD VSS sg13g2_decap_8
XFILLER_10_777 VDD VSS sg13g2_decap_8
XFILLER_108_654 VDD VSS sg13g2_decap_8
XFILLER_30_63 VDD VSS sg13g2_decap_8
XFILLER_107_197 VDD VSS sg13g2_fill_2
XFILLER_107_175 VDD VSS sg13g2_decap_8
XFILLER_107_186 VDD VSS sg13g2_decap_8
XFILLER_2_910 VDD VSS sg13g2_decap_8
XFILLER_111_819 VDD VSS sg13g2_decap_8
XFILLER_1_420 VDD VSS sg13g2_decap_8
XFILLER_2_987 VDD VSS sg13g2_decap_8
XFILLER_1_497 VDD VSS sg13g2_decap_8
XFILLER_7_1036 VDD VSS sg13g2_decap_8
XFILLER_92_703 VDD VSS sg13g2_decap_8
XFILLER_92_714 VDD VSS sg13g2_decap_8
XFILLER_77_788 VDD VSS sg13g2_decap_8
XFILLER_76_254 VDD VSS sg13g2_decap_8
XFILLER_58_980 VDD VSS sg13g2_decap_8
XFILLER_91_213 VDD VSS sg13g2_decap_8
XFILLER_76_298 VDD VSS sg13g2_fill_1
XFILLER_18_833 VDD VSS sg13g2_decap_8
XFILLER_45_641 VDD VSS sg13g2_fill_2
XFILLER_17_343 VDD VSS sg13g2_decap_8
XFILLER_33_847 VDD VSS sg13g2_decap_8
XFILLER_32_357 VDD VSS sg13g2_decap_8
XFILLER_13_560 VDD VSS sg13g2_decap_8
X_2234__285 VDD VSS _2234_/RESET_B sg13g2_tiehi
XFILLER_71_92 VDD VSS sg13g2_fill_2
XFILLER_9_553 VDD VSS sg13g2_decap_8
XFILLER_5_770 VDD VSS sg13g2_decap_8
X_1523_ _1594_/A _1523_/B _1584_/B VDD VSS sg13g2_nor2_1
XFILLER_99_346 VDD VSS sg13g2_decap_8
X_1454_ VSS VDD _1373_/Y _1453_/B _2246_/D _1453_/Y sg13g2_a21oi_1
XFILLER_4_280 VDD VSS sg13g2_decap_8
XFILLER_45_1031 VDD VSS sg13g2_decap_8
XFILLER_68_733 VDD VSS sg13g2_fill_1
XFILLER_68_722 VDD VSS sg13g2_decap_8
XFILLER_110_830 VDD VSS sg13g2_decap_8
XFILLER_56_906 VDD VSS sg13g2_decap_8
X_1385_ _1385_/Y _1385_/A _1465_/C VDD VSS sg13g2_nand2_1
X_2198__144 VDD VSS _2198_/RESET_B sg13g2_tiehi
XFILLER_67_265 VDD VSS sg13g2_decap_4
XFILLER_95_596 VDD VSS sg13g2_decap_8
XFILLER_36_630 VDD VSS sg13g2_decap_8
XFILLER_67_287 VDD VSS sg13g2_decap_8
XFILLER_55_438 VDD VSS sg13g2_decap_8
X_2006_ _2071_/A VDD _2160_/B VSS _2004_/B _2005_/X sg13g2_o21ai_1
XFILLER_82_257 VDD VSS sg13g2_decap_8
XFILLER_64_972 VDD VSS sg13g2_decap_4
XFILLER_35_140 VDD VSS sg13g2_decap_8
XFILLER_91_780 VDD VSS sg13g2_decap_8
XFILLER_51_600 VDD VSS sg13g2_fill_1
XFILLER_24_847 VDD VSS sg13g2_decap_8
XFILLER_63_482 VDD VSS sg13g2_decap_8
XFILLER_51_633 VDD VSS sg13g2_decap_8
XFILLER_23_357 VDD VSS sg13g2_decap_8
XFILLER_50_165 VDD VSS sg13g2_fill_1
XFILLER_13_1008 VDD VSS sg13g2_decap_8
XFILLER_105_602 VDD VSS sg13g2_decap_8
XFILLER_3_707 VDD VSS sg13g2_decap_8
XFILLER_104_112 VDD VSS sg13g2_decap_8
XFILLER_2_217 VDD VSS sg13g2_decap_8
XFILLER_105_679 VDD VSS sg13g2_decap_8
XFILLER_78_508 VDD VSS sg13g2_decap_8
XFILLER_104_167 VDD VSS sg13g2_decap_8
XFILLER_98_390 VDD VSS sg13g2_decap_8
XFILLER_86_563 VDD VSS sg13g2_decap_8
XFILLER_46_416 VDD VSS sg13g2_fill_1
XFILLER_74_736 VDD VSS sg13g2_decap_4
XFILLER_27_630 VDD VSS sg13g2_decap_8
XFILLER_73_257 VDD VSS sg13g2_fill_2
XFILLER_92_14 VDD VSS sg13g2_decap_8
XFILLER_55_950 VDD VSS sg13g2_decap_4
XFILLER_26_140 VDD VSS sg13g2_decap_8
XFILLER_70_920 VDD VSS sg13g2_decap_8
XFILLER_55_994 VDD VSS sg13g2_fill_2
XFILLER_54_460 VDD VSS sg13g2_decap_8
XFILLER_109_1036 VDD VSS sg13g2_decap_8
XFILLER_42_644 VDD VSS sg13g2_decap_8
XFILLER_15_847 VDD VSS sg13g2_decap_8
XFILLER_25_63 VDD VSS sg13g2_decap_8
XFILLER_70_997 VDD VSS sg13g2_decap_8
XFILLER_14_357 VDD VSS sg13g2_decap_8
X_2368__236 VDD VSS _2368_/RESET_B sg13g2_tiehi
XFILLER_109_952 VDD VSS sg13g2_decap_8
XFILLER_10_574 VDD VSS sg13g2_decap_8
XFILLER_41_84 VDD VSS sg13g2_decap_8
XFILLER_6_567 VDD VSS sg13g2_decap_8
XFILLER_29_1015 VDD VSS sg13g2_decap_8
XFILLER_69_508 VDD VSS sg13g2_decap_4
XFILLER_111_616 VDD VSS sg13g2_decap_8
XFILLER_97_839 VDD VSS sg13g2_decap_8
XFILLER_2_784 VDD VSS sg13g2_decap_8
XFILLER_77_530 VDD VSS sg13g2_decap_8
XFILLER_110_126 VDD VSS sg13g2_decap_8
XFILLER_1_294 VDD VSS sg13g2_decap_8
XFILLER_65_703 VDD VSS sg13g2_decap_8
XFILLER_2_56 VDD VSS sg13g2_decap_8
XFILLER_92_533 VDD VSS sg13g2_decap_8
XFILLER_66_70 VDD VSS sg13g2_decap_8
XFILLER_37_427 VDD VSS sg13g2_decap_8
XFILLER_92_544 VDD VSS sg13g2_fill_1
XFILLER_46_961 VDD VSS sg13g2_decap_8
XFILLER_64_268 VDD VSS sg13g2_decap_8
XFILLER_18_630 VDD VSS sg13g2_decap_8
XFILLER_80_739 VDD VSS sg13g2_decap_8
XFILLER_52_419 VDD VSS sg13g2_fill_1
XFILLER_17_140 VDD VSS sg13g2_decap_8
XFILLER_36_1008 VDD VSS sg13g2_decap_8
XFILLER_33_644 VDD VSS sg13g2_decap_8
XFILLER_82_91 VDD VSS sg13g2_decap_8
XFILLER_32_154 VDD VSS sg13g2_decap_8
XFILLER_9_350 VDD VSS sg13g2_decap_8
XFILLER_56_0 VDD VSS sg13g2_decap_8
XFILLER_102_616 VDD VSS sg13g2_decap_8
X_1506_ _1510_/B _1510_/A _1506_/X VDD VSS sg13g2_xor2_1
XFILLER_96_850 VDD VSS sg13g2_decap_8
XFILLER_99_198 VDD VSS sg13g2_decap_8
XFILLER_101_126 VDD VSS sg13g2_decap_8
X_1437_ VDD _2238_/D _1437_/A VSS sg13g2_inv_1
XFILLER_68_530 VDD VSS sg13g2_decap_8
X_1368_ _1368_/Y _1368_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_29_917 VDD VSS sg13g2_decap_8
XFILLER_56_714 VDD VSS sg13g2_decap_8
XFILLER_83_511 VDD VSS sg13g2_decap_8
XFILLER_55_224 VDD VSS sg13g2_decap_8
XFILLER_28_427 VDD VSS sg13g2_decap_8
XFILLER_71_706 VDD VSS sg13g2_decap_8
X_1299_ VDD _2179_/D _1299_/A VSS sg13g2_inv_1
XFILLER_102_35 VDD VSS sg13g2_decap_8
XFILLER_37_994 VDD VSS sg13g2_decap_8
XFILLER_24_644 VDD VSS sg13g2_decap_8
XFILLER_63_290 VDD VSS sg13g2_decap_8
XFILLER_62_28 VDD VSS sg13g2_decap_8
XFILLER_52_997 VDD VSS sg13g2_decap_8
XFILLER_51_463 VDD VSS sg13g2_decap_4
XFILLER_23_154 VDD VSS sg13g2_decap_8
XFILLER_20_861 VDD VSS sg13g2_decap_8
XFILLER_11_21 VDD VSS sg13g2_decap_8
XFILLER_106_944 VDD VSS sg13g2_decap_8
XFILLER_3_504 VDD VSS sg13g2_decap_8
XFILLER_105_421 VDD VSS sg13g2_decap_8
XFILLER_87_14 VDD VSS sg13g2_decap_8
XFILLER_11_98 VDD VSS sg13g2_decap_8
XFILLER_79_828 VDD VSS sg13g2_decap_8
XFILLER_87_850 VDD VSS sg13g2_decap_8
XFILLER_78_349 VDD VSS sg13g2_decap_4
XFILLER_74_500 VDD VSS sg13g2_decap_8
XFILLER_59_574 VDD VSS sg13g2_decap_4
XFILLER_101_671 VDD VSS sg13g2_decap_8
XFILLER_47_736 VDD VSS sg13g2_decap_8
XFILLER_19_427 VDD VSS sg13g2_decap_8
XFILLER_46_213 VDD VSS sg13g2_decap_8
XFILLER_98_1046 VDD VSS sg13g2_decap_8
XFILLER_74_599 VDD VSS sg13g2_decap_8
XFILLER_74_588 VDD VSS sg13g2_decap_8
XFILLER_28_994 VDD VSS sg13g2_decap_8
XFILLER_61_227 VDD VSS sg13g2_decap_8
XFILLER_15_644 VDD VSS sg13g2_decap_8
XFILLER_36_84 VDD VSS sg13g2_decap_8
XFILLER_43_975 VDD VSS sg13g2_decap_8
XFILLER_14_154 VDD VSS sg13g2_decap_8
XFILLER_70_794 VDD VSS sg13g2_decap_8
XFILLER_30_658 VDD VSS sg13g2_decap_8
XFILLER_11_861 VDD VSS sg13g2_decap_8
XFILLER_10_371 VDD VSS sg13g2_decap_8
XFILLER_7_854 VDD VSS sg13g2_decap_8
XFILLER_6_364 VDD VSS sg13g2_decap_8
XFILLER_112_903 VDD VSS sg13g2_decap_8
XFILLER_97_614 VDD VSS sg13g2_decap_8
X_2340_ _2340_/RESET_B VSS VDD _2340_/D _2340_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_111_413 VDD VSS sg13g2_decap_8
XFILLER_69_316 VDD VSS sg13g2_decap_8
XFILLER_97_647 VDD VSS sg13g2_decap_8
XFILLER_42_1001 VDD VSS sg13g2_decap_8
X_2271_ _2271_/RESET_B VSS VDD _2271_/D _2271_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_2_581 VDD VSS sg13g2_decap_8
XFILLER_96_168 VDD VSS sg13g2_decap_8
XFILLER_77_91 VDD VSS sg13g2_decap_8
X_1222_ _2101_/A _1222_/B _1238_/B _1222_/Y VDD VSS sg13g2_nor3_1
XFILLER_65_522 VDD VSS sg13g2_decap_8
XFILLER_37_224 VDD VSS sg13g2_decap_8
XFILLER_38_758 VDD VSS sg13g2_decap_8
XFILLER_19_994 VDD VSS sg13g2_decap_8
XFILLER_52_216 VDD VSS sg13g2_fill_2
XFILLER_92_396 VDD VSS sg13g2_decap_8
XFILLER_34_931 VDD VSS sg13g2_decap_8
XFILLER_45_290 VDD VSS sg13g2_decap_8
XFILLER_61_772 VDD VSS sg13g2_decap_8
XFILLER_33_441 VDD VSS sg13g2_decap_8
XFILLER_61_783 VDD VSS sg13g2_fill_1
X_1986_ VSS VDD _1984_/A _1984_/B _1987_/B _1945_/X sg13g2_a21oi_1
XFILLER_21_658 VDD VSS sg13g2_decap_8
XFILLER_20_168 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_9_clk clkbuf_leaf_9_clk/A _2345_/CLK VDD VSS sg13g2_buf_8
XFILLER_103_903 VDD VSS sg13g2_decap_8
XFILLER_88_614 VDD VSS sg13g2_decap_8
X_2282__175 VDD VSS _2282_/RESET_B sg13g2_tiehi
XFILLER_0_518 VDD VSS sg13g2_decap_8
XFILLER_76_809 VDD VSS sg13g2_decap_8
XFILLER_102_435 VDD VSS sg13g2_decap_8
XFILLER_69_861 VDD VSS sg13g2_decap_8
XFILLER_57_28 VDD VSS sg13g2_fill_1
XFILLER_111_980 VDD VSS sg13g2_decap_8
XFILLER_87_179 VDD VSS sg13g2_decap_4
XFILLER_29_714 VDD VSS sg13g2_decap_8
XFILLER_68_371 VDD VSS sg13g2_fill_1
XFILLER_84_864 VDD VSS sg13g2_decap_8
XFILLER_56_533 VDD VSS sg13g2_decap_4
XFILLER_28_224 VDD VSS sg13g2_decap_8
XFILLER_56_588 VDD VSS sg13g2_decap_8
XFILLER_44_739 VDD VSS sg13g2_decap_8
XFILLER_3_1050 VDD VSS sg13g2_decap_8
XFILLER_83_396 VDD VSS sg13g2_decap_8
XFILLER_71_536 VDD VSS sg13g2_decap_8
XFILLER_73_49 VDD VSS sg13g2_decap_8
XFILLER_25_931 VDD VSS sg13g2_decap_8
XFILLER_37_791 VDD VSS sg13g2_decap_8
XFILLER_58_1052 VDD VSS sg13g2_decap_8
XFILLER_52_772 VDD VSS sg13g2_decap_8
XFILLER_19_1036 VDD VSS sg13g2_decap_8
XFILLER_24_441 VDD VSS sg13g2_decap_8
XFILLER_106_1028 VDD VSS sg13g2_decap_8
XFILLER_40_956 VDD VSS sg13g2_decap_8
XFILLER_12_658 VDD VSS sg13g2_decap_8
XFILLER_11_168 VDD VSS sg13g2_decap_8
XFILLER_22_42 VDD VSS sg13g2_decap_8
XFILLER_98_35 VDD VSS sg13g2_decap_8
XFILLER_3_301 VDD VSS sg13g2_decap_8
XFILLER_106_741 VDD VSS sg13g2_decap_8
XFILLER_65_1001 VDD VSS sg13g2_decap_8
XFILLER_4_868 VDD VSS sg13g2_decap_8
XFILLER_3_378 VDD VSS sg13g2_decap_8
XFILLER_26_1029 VDD VSS sg13g2_decap_8
XFILLER_66_308 VDD VSS sg13g2_decap_8
XFILLER_93_105 VDD VSS sg13g2_decap_8
XFILLER_101_490 VDD VSS sg13g2_fill_1
XFILLER_19_224 VDD VSS sg13g2_decap_8
XFILLER_75_897 VDD VSS sg13g2_decap_8
XFILLER_74_352 VDD VSS sg13g2_decap_8
XFILLER_35_728 VDD VSS sg13g2_decap_8
XFILLER_74_396 VDD VSS sg13g2_fill_1
XFILLER_62_547 VDD VSS sg13g2_decap_8
XFILLER_28_791 VDD VSS sg13g2_decap_8
XFILLER_16_931 VDD VSS sg13g2_decap_8
XFILLER_34_238 VDD VSS sg13g2_decap_8
XFILLER_43_772 VDD VSS sg13g2_decap_8
XFILLER_15_441 VDD VSS sg13g2_decap_8
XFILLER_70_591 VDD VSS sg13g2_decap_8
XFILLER_97_7 VDD VSS sg13g2_decap_8
XFILLER_31_945 VDD VSS sg13g2_decap_8
X_1840_ _1934_/A _2244_/Q _2203_/Q VDD VSS sg13g2_nand2b_1
X_2228__84 VDD VSS _2228__84/L_HI sg13g2_tiehi
XFILLER_30_455 VDD VSS sg13g2_decap_8
X_1771_ _1770_/A VDD _1877_/A VSS _1888_/A _1770_/B sg13g2_o21ai_1
XFILLER_8_77 VDD VSS sg13g2_decap_8
XFILLER_7_651 VDD VSS sg13g2_decap_8
XFILLER_6_161 VDD VSS sg13g2_decap_8
XFILLER_112_700 VDD VSS sg13g2_decap_8
XFILLER_97_400 VDD VSS sg13g2_decap_8
XFILLER_98_945 VDD VSS sg13g2_decap_4
X_2323_ _2323_/RESET_B VSS VDD _2323_/D _2323_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_111_210 VDD VSS sg13g2_decap_8
XFILLER_69_113 VDD VSS sg13g2_decap_8
XFILLER_112_777 VDD VSS sg13g2_decap_8
XFILLER_85_617 VDD VSS sg13g2_decap_8
XFILLER_97_466 VDD VSS sg13g2_decap_8
XFILLER_58_809 VDD VSS sg13g2_decap_8
XFILLER_111_287 VDD VSS sg13g2_decap_8
XFILLER_97_499 VDD VSS sg13g2_decap_8
XFILLER_97_488 VDD VSS sg13g2_decap_4
XFILLER_84_105 VDD VSS sg13g2_decap_8
X_2254_ _2254_/RESET_B VSS VDD _2254_/D _2254_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_66_831 VDD VSS sg13g2_decap_8
XFILLER_84_149 VDD VSS sg13g2_decap_8
XFILLER_66_842 VDD VSS sg13g2_fill_2
X_2185_ _2185_/RESET_B VSS VDD _2185_/D _2185_/Q clkload8/A sg13g2_dfrbpq_1
X_1205_ VDD _2110_/A _1510_/A VSS sg13g2_inv_1
XFILLER_38_555 VDD VSS sg13g2_decap_8
XFILLER_19_0 VDD VSS sg13g2_decap_8
XFILLER_93_672 VDD VSS sg13g2_decap_8
XFILLER_26_728 VDD VSS sg13g2_decap_8
XFILLER_81_856 VDD VSS sg13g2_fill_1
XFILLER_92_171 VDD VSS sg13g2_decap_8
XFILLER_65_385 VDD VSS sg13g2_decap_8
XFILLER_19_791 VDD VSS sg13g2_decap_8
XFILLER_25_238 VDD VSS sg13g2_decap_8
XFILLER_80_355 VDD VSS sg13g2_decap_8
XFILLER_22_945 VDD VSS sg13g2_decap_8
XFILLER_21_455 VDD VSS sg13g2_decap_8
XFILLER_105_1050 VDD VSS sg13g2_decap_8
X_1969_ _1968_/Y VDD _1973_/B VSS _1966_/A _1966_/B sg13g2_o21ai_1
XFILLER_107_527 VDD VSS sg13g2_decap_8
XFILLER_103_711 VDD VSS sg13g2_fill_2
XFILLER_89_901 VDD VSS sg13g2_decap_8
XFILLER_108_56 VDD VSS sg13g2_decap_8
XFILLER_1_805 VDD VSS sg13g2_decap_8
XFILLER_88_422 VDD VSS sg13g2_decap_8
XFILLER_0_315 VDD VSS sg13g2_decap_8
XFILLER_68_49 VDD VSS sg13g2_decap_8
XFILLER_89_989 VDD VSS sg13g2_decap_8
XFILLER_103_777 VDD VSS sg13g2_decap_8
XFILLER_76_617 VDD VSS sg13g2_decap_4
XFILLER_102_276 VDD VSS sg13g2_decap_8
XFILLER_102_287 VDD VSS sg13g2_decap_8
XFILLER_75_105 VDD VSS sg13g2_decap_8
XFILLER_29_511 VDD VSS sg13g2_decap_8
XFILLER_112_1043 VDD VSS sg13g2_decap_8
XFILLER_91_609 VDD VSS sg13g2_decap_8
XFILLER_68_190 VDD VSS sg13g2_decap_8
XFILLER_84_683 VDD VSS sg13g2_decap_8
XFILLER_72_801 VDD VSS sg13g2_decap_8
XFILLER_29_588 VDD VSS sg13g2_decap_8
XFILLER_56_363 VDD VSS sg13g2_decap_8
XFILLER_17_728 VDD VSS sg13g2_decap_8
XFILLER_71_322 VDD VSS sg13g2_fill_2
XFILLER_16_238 VDD VSS sg13g2_decap_8
XFILLER_17_42 VDD VSS sg13g2_decap_8
XFILLER_44_536 VDD VSS sg13g2_decap_8
X_2371__265 VDD VSS _2371_/RESET_B sg13g2_tiehi
XIO_BOND_in_data_pads\[4\].in_data_pad in_data_PADs[4] bondpad_70x70
XFILLER_13_945 VDD VSS sg13g2_decap_8
XFILLER_40_753 VDD VSS sg13g2_decap_8
XFILLER_12_455 VDD VSS sg13g2_decap_8
XFILLER_32_1022 VDD VSS sg13g2_decap_8
XFILLER_9_938 VDD VSS sg13g2_decap_8
XFILLER_33_63 VDD VSS sg13g2_decap_8
XFILLER_8_448 VDD VSS sg13g2_decap_8
XFILLER_4_665 VDD VSS sg13g2_decap_8
XFILLER_79_433 VDD VSS sg13g2_decap_8
XFILLER_3_175 VDD VSS sg13g2_decap_8
XFILLER_95_959 VDD VSS sg13g2_decap_8
XFILLER_67_628 VDD VSS sg13g2_decap_8
XFILLER_0_882 VDD VSS sg13g2_decap_8
XFILLER_66_105 VDD VSS sg13g2_decap_8
XFILLER_94_447 VDD VSS sg13g2_decap_8
XFILLER_48_842 VDD VSS sg13g2_decap_4
XFILLER_12_7 VDD VSS sg13g2_decap_8
XFILLER_58_93 VDD VSS sg13g2_decap_8
XFILLER_75_672 VDD VSS sg13g2_decap_8
XFILLER_81_119 VDD VSS sg13g2_fill_2
XFILLER_47_352 VDD VSS sg13g2_decap_4
XFILLER_74_70 VDD VSS sg13g2_decap_8
XFILLER_35_525 VDD VSS sg13g2_decap_8
XFILLER_47_385 VDD VSS sg13g2_decap_8
XFILLER_90_675 VDD VSS sg13g2_decap_8
XFILLER_63_867 VDD VSS sg13g2_decap_8
XFILLER_62_366 VDD VSS sg13g2_fill_1
XFILLER_62_344 VDD VSS sg13g2_decap_8
XFILLER_50_539 VDD VSS sg13g2_decap_8
XFILLER_31_742 VDD VSS sg13g2_decap_8
XFILLER_90_91 VDD VSS sg13g2_decap_8
XFILLER_30_252 VDD VSS sg13g2_decap_8
X_1823_ _1823_/B _1823_/A _1878_/B VDD VSS sg13g2_xor2_1
X_1754_ VSS VDD _1750_/A _1752_/Y _1754_/Y _1753_/Y sg13g2_a21oi_1
Xhold426 _2240_/Q VDD VSS hold426/X sg13g2_dlygate4sd3_1
Xhold404 _2195_/Q VDD VSS hold404/X sg13g2_dlygate4sd3_1
Xhold415 _2361_/Q VDD VSS _1500_/B sg13g2_dlygate4sd3_1
Xhold448 _2230_/Q VDD VSS _1418_/A sg13g2_dlygate4sd3_1
X_1685_ _1685_/B _2313_/Q _1686_/B VDD VSS sg13g2_xor2_1
Xhold437 _2300_/Q VDD VSS hold437/X sg13g2_dlygate4sd3_1
Xhold459 _2250_/Q VDD VSS _1461_/A sg13g2_dlygate4sd3_1
XFILLER_48_1051 VDD VSS sg13g2_decap_8
XFILLER_100_703 VDD VSS sg13g2_decap_8
XFILLER_86_937 VDD VSS sg13g2_decap_8
XFILLER_112_574 VDD VSS sg13g2_decap_8
XFILLER_97_263 VDD VSS sg13g2_decap_8
X_2306_ _2306__87/L_HI VSS VDD _2306_/D _2306_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_85_447 VDD VSS sg13g2_decap_8
X_2237_ _2237_/RESET_B VSS VDD _2237_/D _2237_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_72_119 VDD VSS sg13g2_fill_1
XFILLER_54_801 VDD VSS sg13g2_decap_8
XFILLER_39_864 VDD VSS sg13g2_decap_8
XFILLER_38_341 VDD VSS sg13g2_decap_8
X_2168_ _2168_/RESET_B VSS VDD _2168_/D _2168_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_26_525 VDD VSS sg13g2_decap_8
XFILLER_54_878 VDD VSS sg13g2_decap_8
X_2099_ _2099_/B _2099_/A _2099_/X VDD VSS sg13g2_xor2_1
XFILLER_80_185 VDD VSS sg13g2_decap_8
XFILLER_110_35 VDD VSS sg13g2_decap_8
XFILLER_22_742 VDD VSS sg13g2_decap_8
XFILLER_70_28 VDD VSS sg13g2_decap_8
XFILLER_21_252 VDD VSS sg13g2_decap_8
XFILLER_10_959 VDD VSS sg13g2_decap_8
XFILLER_108_836 VDD VSS sg13g2_decap_8
XFILLER_107_346 VDD VSS sg13g2_decap_8
XFILLER_1_602 VDD VSS sg13g2_decap_8
XFILLER_0_112 VDD VSS sg13g2_decap_8
XFILLER_95_14 VDD VSS sg13g2_decap_8
XFILLER_77_926 VDD VSS sg13g2_decap_8
XFILLER_103_574 VDD VSS sg13g2_decap_8
XFILLER_62_1059 VDD VSS sg13g2_fill_2
XFILLER_1_679 VDD VSS sg13g2_decap_8
XFILLER_0_189 VDD VSS sg13g2_decap_8
XFILLER_76_469 VDD VSS sg13g2_decap_8
XFILLER_28_63 VDD VSS sg13g2_decap_8
XFILLER_17_525 VDD VSS sg13g2_decap_8
XFILLER_29_385 VDD VSS sg13g2_decap_8
XFILLER_44_322 VDD VSS sg13g2_decap_8
XFILLER_72_675 VDD VSS sg13g2_decap_8
XFILLER_45_889 VDD VSS sg13g2_fill_2
XFILLER_32_539 VDD VSS sg13g2_decap_8
XFILLER_44_399 VDD VSS sg13g2_decap_4
XFILLER_13_742 VDD VSS sg13g2_decap_8
XFILLER_44_84 VDD VSS sg13g2_decap_8
XFILLER_40_550 VDD VSS sg13g2_decap_8
XFILLER_12_252 VDD VSS sg13g2_decap_8
XFILLER_9_735 VDD VSS sg13g2_decap_8
XFILLER_8_245 VDD VSS sg13g2_decap_8
XFILLER_60_94 VDD VSS sg13g2_decap_4
XFILLER_5_952 VDD VSS sg13g2_decap_8
XFILLER_107_891 VDD VSS sg13g2_decap_8
X_1470_ _1367_/A VDD _1470_/Y VSS _1373_/A _1479_/A2 sg13g2_o21ai_1
X_2343__131 VDD VSS _2343_/RESET_B sg13g2_tiehi
XFILLER_4_462 VDD VSS sg13g2_decap_8
XFILLER_5_56 VDD VSS sg13g2_decap_8
XFILLER_69_92 VDD VSS sg13g2_decap_8
XFILLER_68_904 VDD VSS sg13g2_decap_8
XFILLER_39_105 VDD VSS sg13g2_decap_8
XFILLER_67_436 VDD VSS sg13g2_decap_8
XFILLER_76_970 VDD VSS sg13g2_decap_8
XFILLER_36_812 VDD VSS sg13g2_decap_8
XFILLER_91_940 VDD VSS sg13g2_decap_8
X_2022_ _2009_/X _2021_/X _2022_/S _2022_/X VDD VSS sg13g2_mux2_1
XFILLER_85_91 VDD VSS sg13g2_decap_8
XFILLER_48_694 VDD VSS sg13g2_decap_8
XFILLER_35_322 VDD VSS sg13g2_decap_8
XFILLER_90_450 VDD VSS sg13g2_decap_8
XFILLER_63_642 VDD VSS sg13g2_decap_8
XFILLER_36_889 VDD VSS sg13g2_decap_8
XFILLER_62_141 VDD VSS sg13g2_decap_8
XFILLER_90_483 VDD VSS sg13g2_decap_8
XFILLER_39_1039 VDD VSS sg13g2_decap_8
XFILLER_23_539 VDD VSS sg13g2_decap_8
XFILLER_35_399 VDD VSS sg13g2_decap_8
XFILLER_62_185 VDD VSS sg13g2_decap_8
XFILLER_50_325 VDD VSS sg13g2_decap_8
XFILLER_86_0 VDD VSS sg13g2_decap_8
XFILLER_102_1020 VDD VSS sg13g2_decap_8
X_1806_ _1812_/A _1812_/B _1806_/Y VDD VSS sg13g2_nor2_1
XFILLER_15_1050 VDD VSS sg13g2_decap_8
X_1737_ _1915_/B _2230_/Q _2238_/Q VDD VSS sg13g2_xnor2_1
X_1668_ _1674_/B _2335_/Q _2327_/Q _2350_/Q _2342_/Q _1677_/A _1668_/X VDD VSS sg13g2_mux4_1
XFILLER_104_349 VDD VSS sg13g2_decap_8
XFILLER_59_915 VDD VSS sg13g2_decap_8
XFILLER_112_371 VDD VSS sg13g2_decap_8
X_1599_ _2275_/Q _2290_/Q _1600_/B VDD VSS sg13g2_xor2_1
XFILLER_86_767 VDD VSS sg13g2_decap_8
XFILLER_105_35 VDD VSS sg13g2_decap_8
XFILLER_58_436 VDD VSS sg13g2_decap_8
XFILLER_85_266 VDD VSS sg13g2_decap_8
XFILLER_22_1043 VDD VSS sg13g2_decap_8
XFILLER_39_661 VDD VSS sg13g2_decap_8
XFILLER_27_812 VDD VSS sg13g2_decap_8
XFILLER_65_28 VDD VSS sg13g2_decap_8
XFILLER_100_588 VDD VSS sg13g2_decap_8
XFILLER_85_299 VDD VSS sg13g2_decap_8
XFILLER_73_428 VDD VSS sg13g2_decap_8
XFILLER_67_992 VDD VSS sg13g2_decap_8
XFILLER_26_322 VDD VSS sg13g2_decap_8
XFILLER_38_182 VDD VSS sg13g2_decap_8
XFILLER_81_461 VDD VSS sg13g2_decap_8
XFILLER_42_826 VDD VSS sg13g2_decap_8
XFILLER_27_889 VDD VSS sg13g2_decap_8
XFILLER_14_539 VDD VSS sg13g2_decap_8
XFILLER_81_49 VDD VSS sg13g2_decap_8
XFILLER_53_196 VDD VSS sg13g2_decap_8
XFILLER_26_399 VDD VSS sg13g2_decap_8
XFILLER_41_336 VDD VSS sg13g2_decap_8
XFILLER_14_21 VDD VSS sg13g2_decap_8
XFILLER_14_98 VDD VSS sg13g2_decap_8
XFILLER_10_756 VDD VSS sg13g2_decap_8
XFILLER_108_633 VDD VSS sg13g2_decap_8
XFILLER_6_749 VDD VSS sg13g2_decap_8
XFILLER_107_154 VDD VSS sg13g2_decap_8
XFILLER_5_259 VDD VSS sg13g2_decap_8
XFILLER_30_42 VDD VSS sg13g2_decap_8
XFILLER_2_966 VDD VSS sg13g2_decap_8
XFILLER_104_872 VDD VSS sg13g2_fill_2
XFILLER_89_572 VDD VSS sg13g2_decap_4
XFILLER_77_723 VDD VSS sg13g2_decap_4
XFILLER_110_308 VDD VSS sg13g2_fill_2
XFILLER_110_319 VDD VSS sg13g2_decap_8
XFILLER_1_476 VDD VSS sg13g2_decap_8
XFILLER_7_1015 VDD VSS sg13g2_decap_8
XFILLER_77_767 VDD VSS sg13g2_decap_8
XFILLER_76_233 VDD VSS sg13g2_decap_8
XFILLER_39_84 VDD VSS sg13g2_decap_8
XFILLER_49_447 VDD VSS sg13g2_decap_8
XFILLER_37_609 VDD VSS sg13g2_decap_8
XFILLER_18_812 VDD VSS sg13g2_decap_8
XFILLER_45_631 VDD VSS sg13g2_fill_1
XFILLER_17_322 VDD VSS sg13g2_decap_8
XFILLER_36_119 VDD VSS sg13g2_decap_8
XFILLER_91_269 VDD VSS sg13g2_decap_8
XFILLER_44_141 VDD VSS sg13g2_decap_8
XFILLER_29_182 VDD VSS sg13g2_decap_8
XFILLER_72_483 VDD VSS sg13g2_decap_8
XFILLER_60_623 VDD VSS sg13g2_fill_2
XFILLER_60_612 VDD VSS sg13g2_decap_8
XFILLER_45_697 VDD VSS sg13g2_decap_8
XFILLER_33_826 VDD VSS sg13g2_decap_8
XFILLER_18_889 VDD VSS sg13g2_decap_8
XFILLER_17_399 VDD VSS sg13g2_decap_8
XFILLER_32_336 VDD VSS sg13g2_decap_8
XFILLER_41_881 VDD VSS sg13g2_decap_8
XFILLER_9_532 VDD VSS sg13g2_decap_8
XFILLER_40_391 VDD VSS sg13g2_decap_8
XFILLER_99_325 VDD VSS sg13g2_decap_8
X_1522_ _1522_/Y _1592_/A _1589_/B VDD VSS sg13g2_nand2b_1
X_1453_ _1453_/A _1453_/B _1453_/Y VDD VSS sg13g2_nor2_1
XFILLER_45_1010 VDD VSS sg13g2_decap_8
XFILLER_68_701 VDD VSS sg13g2_decap_8
X_1384_ _1383_/Y VDD _2216_/D VSS _1367_/B _1382_/Y sg13g2_o21ai_1
XFILLER_110_886 VDD VSS sg13g2_decap_8
XFILLER_95_575 VDD VSS sg13g2_decap_8
XFILLER_68_789 VDD VSS sg13g2_fill_2
XFILLER_68_778 VDD VSS sg13g2_decap_8
XFILLER_28_609 VDD VSS sg13g2_decap_8
XFILLER_67_244 VDD VSS sg13g2_decap_8
XFILLER_55_406 VDD VSS sg13g2_fill_2
XFILLER_83_726 VDD VSS sg13g2_decap_8
XFILLER_49_981 VDD VSS sg13g2_decap_8
XFILLER_55_417 VDD VSS sg13g2_decap_8
XFILLER_27_119 VDD VSS sg13g2_decap_8
X_2005_ _2071_/B _2005_/B _2005_/C _2005_/D _2005_/X VDD VSS sg13g2_or4_1
XFILLER_82_236 VDD VSS sg13g2_decap_8
XFILLER_64_951 VDD VSS sg13g2_decap_8
X_2278__191 VDD VSS _2278_/RESET_B sg13g2_tiehi
XFILLER_51_612 VDD VSS sg13g2_decap_8
XFILLER_36_686 VDD VSS sg13g2_decap_8
XFILLER_24_826 VDD VSS sg13g2_decap_8
XFILLER_63_461 VDD VSS sg13g2_decap_8
XFILLER_23_336 VDD VSS sg13g2_decap_8
XFILLER_35_196 VDD VSS sg13g2_decap_8
XFILLER_51_689 VDD VSS sg13g2_decap_8
XFILLER_50_144 VDD VSS sg13g2_decap_8
XFILLER_50_188 VDD VSS sg13g2_decap_8
XFILLER_105_658 VDD VSS sg13g2_decap_8
XFILLER_101_842 VDD VSS sg13g2_fill_2
XFILLER_86_542 VDD VSS sg13g2_decap_8
XFILLER_86_531 VDD VSS sg13g2_decap_4
XFILLER_76_49 VDD VSS sg13g2_decap_8
XFILLER_58_222 VDD VSS sg13g2_fill_2
XFILLER_47_929 VDD VSS sg13g2_fill_2
XFILLER_59_789 VDD VSS sg13g2_decap_8
XFILLER_19_609 VDD VSS sg13g2_decap_8
XFILLER_100_396 VDD VSS sg13g2_fill_2
XFILLER_100_363 VDD VSS sg13g2_decap_8
XFILLER_58_288 VDD VSS sg13g2_decap_8
XFILLER_18_119 VDD VSS sg13g2_decap_8
XFILLER_73_236 VDD VSS sg13g2_decap_8
XFILLER_55_973 VDD VSS sg13g2_decap_8
XFILLER_27_686 VDD VSS sg13g2_decap_8
XFILLER_15_826 VDD VSS sg13g2_decap_8
XFILLER_109_1015 VDD VSS sg13g2_decap_8
XFILLER_82_792 VDD VSS sg13g2_decap_8
XFILLER_81_291 VDD VSS sg13g2_decap_8
XFILLER_42_623 VDD VSS sg13g2_decap_8
XFILLER_14_336 VDD VSS sg13g2_decap_8
XFILLER_25_42 VDD VSS sg13g2_decap_8
XFILLER_26_196 VDD VSS sg13g2_decap_8
XFILLER_70_976 VDD VSS sg13g2_decap_8
XFILLER_41_133 VDD VSS sg13g2_decap_8
XFILLER_41_188 VDD VSS sg13g2_decap_8
XFILLER_10_553 VDD VSS sg13g2_decap_8
XFILLER_109_931 VDD VSS sg13g2_decap_8
XFILLER_41_63 VDD VSS sg13g2_decap_8
XFILLER_6_546 VDD VSS sg13g2_decap_8
XFILLER_108_485 VDD VSS sg13g2_decap_8
XFILLER_68_1054 VDD VSS sg13g2_decap_8
XFILLER_110_105 VDD VSS sg13g2_decap_8
XFILLER_2_763 VDD VSS sg13g2_decap_8
X_2301__107 VDD VSS _2301_/RESET_B sg13g2_tiehi
XFILLER_89_391 VDD VSS sg13g2_decap_8
XFILLER_1_273 VDD VSS sg13g2_decap_8
XFILLER_2_35 VDD VSS sg13g2_decap_8
XFILLER_37_406 VDD VSS sg13g2_decap_8
XFILLER_77_586 VDD VSS sg13g2_decap_8
XFILLER_92_512 VDD VSS sg13g2_decap_8
X_2352__89 VDD VSS _2352__89/L_HI sg13g2_tiehi
XFILLER_49_288 VDD VSS sg13g2_decap_8
XFILLER_65_759 VDD VSS sg13g2_decap_8
XFILLER_64_247 VDD VSS sg13g2_decap_8
XFILLER_75_1003 VDD VSS sg13g2_decap_8
XFILLER_18_686 VDD VSS sg13g2_decap_8
XFILLER_33_623 VDD VSS sg13g2_decap_8
XFILLER_17_196 VDD VSS sg13g2_decap_8
XFILLER_45_483 VDD VSS sg13g2_decap_8
XFILLER_82_70 VDD VSS sg13g2_decap_8
XFILLER_61_965 VDD VSS sg13g2_decap_4
XFILLER_60_442 VDD VSS sg13g2_decap_8
XFILLER_32_133 VDD VSS sg13g2_decap_8
XFILLER_99_133 VDD VSS sg13g2_decap_8
X_1505_ VSS VDD _2110_/A _1514_/A _2269_/D _1504_/Y sg13g2_a21oi_1
XFILLER_49_0 VDD VSS sg13g2_decap_8
XFILLER_99_177 VDD VSS sg13g2_decap_8
XFILLER_101_105 VDD VSS sg13g2_decap_8
X_1436_ _1437_/A _1429_/Y hold477/X _1429_/B _1376_/A VDD VSS sg13g2_a22oi_1
X_1367_ _1367_/A _1367_/B _1389_/B VDD VSS sg13g2_and2_1
XFILLER_28_406 VDD VSS sg13g2_decap_8
XFILLER_110_683 VDD VSS sg13g2_decap_8
XFILLER_68_586 VDD VSS sg13g2_decap_8
XFILLER_55_203 VDD VSS sg13g2_decap_8
X_1298_ _1298_/Y _1482_/B1 hold320/X _1482_/A2 _2343_/Q VDD VSS sg13g2_a22oi_1
XFILLER_83_578 VDD VSS sg13g2_decap_8
XFILLER_102_14 VDD VSS sg13g2_decap_8
XFILLER_37_973 VDD VSS sg13g2_decap_8
XFILLER_64_781 VDD VSS sg13g2_decap_8
XFILLER_52_943 VDD VSS sg13g2_decap_8
XFILLER_24_623 VDD VSS sg13g2_decap_8
XFILLER_36_483 VDD VSS sg13g2_decap_8
XFILLER_52_976 VDD VSS sg13g2_decap_8
XFILLER_52_965 VDD VSS sg13g2_fill_2
XFILLER_23_133 VDD VSS sg13g2_decap_8
XFILLER_20_840 VDD VSS sg13g2_decap_8
XFILLER_106_923 VDD VSS sg13g2_decap_8
XFILLER_105_400 VDD VSS sg13g2_decap_8
XFILLER_11_77 VDD VSS sg13g2_decap_8
XFILLER_105_499 VDD VSS sg13g2_fill_1
XFILLER_78_328 VDD VSS sg13g2_decap_8
XFILLER_59_553 VDD VSS sg13g2_decap_8
XFILLER_98_1025 VDD VSS sg13g2_decap_8
XFILLER_101_661 VDD VSS sg13g2_fill_1
XFILLER_47_726 VDD VSS sg13g2_decap_4
XFILLER_19_406 VDD VSS sg13g2_decap_8
XFILLER_4_1029 VDD VSS sg13g2_decap_8
XFILLER_74_567 VDD VSS sg13g2_decap_8
XFILLER_28_973 VDD VSS sg13g2_decap_8
XFILLER_61_206 VDD VSS sg13g2_decap_8
XFILLER_36_63 VDD VSS sg13g2_decap_8
XFILLER_43_954 VDD VSS sg13g2_decap_8
XFILLER_15_623 VDD VSS sg13g2_decap_8
XFILLER_27_483 VDD VSS sg13g2_decap_8
XFILLER_70_773 VDD VSS sg13g2_decap_8
XFILLER_14_133 VDD VSS sg13g2_decap_8
XFILLER_30_637 VDD VSS sg13g2_decap_8
XFILLER_52_40 VDD VSS sg13g2_decap_8
XFILLER_42_475 VDD VSS sg13g2_decap_4
XFILLER_11_840 VDD VSS sg13g2_decap_8
XFILLER_52_62 VDD VSS sg13g2_decap_8
XFILLER_10_350 VDD VSS sg13g2_decap_8
XFILLER_7_833 VDD VSS sg13g2_decap_8
XFILLER_6_343 VDD VSS sg13g2_decap_8
XFILLER_108_271 VDD VSS sg13g2_decap_8
XFILLER_2_560 VDD VSS sg13g2_decap_8
XFILLER_42_7 VDD VSS sg13g2_decap_8
XFILLER_112_959 VDD VSS sg13g2_decap_8
X_2270_ _2270_/RESET_B VSS VDD _2270_/D _2270_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_111_469 VDD VSS sg13g2_decap_8
XFILLER_96_147 VDD VSS sg13g2_decap_8
XFILLER_77_70 VDD VSS sg13g2_decap_8
X_1221_ _1238_/B _2102_/A _1221_/B VDD VSS sg13g2_nand2_1
XFILLER_93_832 VDD VSS sg13g2_decap_8
XFILLER_78_895 VDD VSS sg13g2_decap_8
XFILLER_42_1057 VDD VSS sg13g2_decap_4
XFILLER_38_737 VDD VSS sg13g2_decap_8
XFILLER_65_501 VDD VSS sg13g2_decap_8
XFILLER_37_203 VDD VSS sg13g2_decap_8
XFILLER_92_375 VDD VSS sg13g2_decap_8
XFILLER_53_718 VDD VSS sg13g2_decap_8
XFILLER_53_729 VDD VSS sg13g2_fill_2
XFILLER_34_910 VDD VSS sg13g2_decap_8
XFILLER_19_973 VDD VSS sg13g2_decap_8
XFILLER_80_537 VDD VSS sg13g2_decap_8
XFILLER_93_91 VDD VSS sg13g2_decap_8
XFILLER_18_483 VDD VSS sg13g2_decap_8
XFILLER_33_420 VDD VSS sg13g2_decap_8
XFILLER_34_987 VDD VSS sg13g2_decap_8
XFILLER_21_637 VDD VSS sg13g2_decap_8
XFILLER_33_497 VDD VSS sg13g2_decap_8
X_1985_ _1987_/A _1985_/A _1985_/B VDD VSS sg13g2_xnor2_1
XFILLER_20_147 VDD VSS sg13g2_decap_8
X_2167__206 VDD VSS _2167_/RESET_B sg13g2_tiehi
XFILLER_107_709 VDD VSS sg13g2_decap_8
X_2247__252 VDD VSS _2247_/RESET_B sg13g2_tiehi
XFILLER_102_403 VDD VSS sg13g2_decap_8
XFILLER_103_959 VDD VSS sg13g2_decap_8
XFILLER_87_125 VDD VSS sg13g2_fill_1
XIO_BOND_clk_pad clk_PAD bondpad_70x70
X_1419_ _1418_/Y VDD _2230_/D VSS _1376_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_87_158 VDD VSS sg13g2_decap_8
XFILLER_68_361 VDD VSS sg13g2_fill_2
XFILLER_56_512 VDD VSS sg13g2_decap_8
XFILLER_28_203 VDD VSS sg13g2_decap_8
XFILLER_110_480 VDD VSS sg13g2_decap_8
XFILLER_83_353 VDD VSS sg13g2_fill_1
XFILLER_73_28 VDD VSS sg13g2_decap_8
XFILLER_56_567 VDD VSS sg13g2_decap_8
XFILLER_44_718 VDD VSS sg13g2_decap_8
XFILLER_37_770 VDD VSS sg13g2_decap_8
XFILLER_25_910 VDD VSS sg13g2_decap_8
XFILLER_24_420 VDD VSS sg13g2_decap_8
XFILLER_36_280 VDD VSS sg13g2_decap_8
XFILLER_43_217 VDD VSS sg13g2_decap_8
XFILLER_43_228 VDD VSS sg13g2_fill_2
XFILLER_25_987 VDD VSS sg13g2_decap_8
XFILLER_52_751 VDD VSS sg13g2_decap_8
XFILLER_19_1015 VDD VSS sg13g2_decap_8
XFILLER_106_1007 VDD VSS sg13g2_decap_8
XFILLER_40_935 VDD VSS sg13g2_decap_8
XFILLER_12_637 VDD VSS sg13g2_decap_8
XFILLER_24_497 VDD VSS sg13g2_decap_8
XFILLER_11_147 VDD VSS sg13g2_decap_8
XFILLER_22_21 VDD VSS sg13g2_decap_8
XFILLER_98_14 VDD VSS sg13g2_decap_8
XFILLER_22_98 VDD VSS sg13g2_decap_8
XFILLER_106_720 VDD VSS sg13g2_decap_8
XFILLER_4_847 VDD VSS sg13g2_decap_8
XFILLER_3_357 VDD VSS sg13g2_decap_8
XFILLER_106_797 VDD VSS sg13g2_decap_8
XFILLER_105_263 VDD VSS sg13g2_decap_8
XFILLER_65_1057 VDD VSS sg13g2_decap_4
XFILLER_26_1008 VDD VSS sg13g2_decap_8
XFILLER_78_147 VDD VSS sg13g2_decap_8
XFILLER_78_158 VDD VSS sg13g2_fill_2
XFILLER_102_970 VDD VSS sg13g2_decap_8
XFILLER_94_629 VDD VSS sg13g2_decap_8
XFILLER_59_383 VDD VSS sg13g2_decap_8
XFILLER_19_203 VDD VSS sg13g2_decap_8
XFILLER_47_545 VDD VSS sg13g2_decap_8
XFILLER_90_813 VDD VSS sg13g2_decap_8
XFILLER_75_876 VDD VSS sg13g2_decap_8
XFILLER_35_707 VDD VSS sg13g2_decap_8
XFILLER_28_770 VDD VSS sg13g2_decap_8
XFILLER_16_910 VDD VSS sg13g2_decap_8
XFILLER_47_84 VDD VSS sg13g2_decap_8
XFILLER_62_526 VDD VSS sg13g2_decap_8
XFILLER_15_420 VDD VSS sg13g2_decap_8
XFILLER_27_280 VDD VSS sg13g2_decap_8
XFILLER_34_217 VDD VSS sg13g2_decap_8
XFILLER_43_751 VDD VSS sg13g2_decap_8
XFILLER_16_987 VDD VSS sg13g2_decap_8
XFILLER_72_1039 VDD VSS sg13g2_decap_8
XFILLER_70_570 VDD VSS sg13g2_decap_8
XFILLER_31_924 VDD VSS sg13g2_decap_8
XFILLER_63_83 VDD VSS sg13g2_decap_8
XFILLER_15_497 VDD VSS sg13g2_decap_8
XFILLER_30_434 VDD VSS sg13g2_decap_8
XFILLER_42_294 VDD VSS sg13g2_decap_8
X_1770_ _1888_/B _1770_/A _1770_/B VDD VSS sg13g2_nand2_1
XFILLER_8_56 VDD VSS sg13g2_decap_8
XFILLER_7_630 VDD VSS sg13g2_decap_8
XFILLER_6_140 VDD VSS sg13g2_decap_8
XFILLER_98_924 VDD VSS sg13g2_decap_8
X_2322_ _2322_/RESET_B VSS VDD _2322_/D _2322_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_88_91 VDD VSS sg13g2_decap_8
XFILLER_112_756 VDD VSS sg13g2_decap_8
XFILLER_97_445 VDD VSS sg13g2_decap_8
XFILLER_111_266 VDD VSS sg13g2_decap_8
XFILLER_84_128 VDD VSS sg13g2_fill_1
X_2253_ _2253_/RESET_B VSS VDD _2253_/D _2253_/Q clkload0/A sg13g2_dfrbpq_1
XFILLER_66_810 VDD VSS sg13g2_decap_8
X_2184_ _2184_/RESET_B VSS VDD _2184_/D _2184_/Q _2372_/CLK sg13g2_dfrbpq_1
X_1204_ VDD _1204_/Y _2309_/Q VSS sg13g2_inv_1
XFILLER_65_320 VDD VSS sg13g2_decap_8
XFILLER_26_707 VDD VSS sg13g2_decap_8
XFILLER_65_364 VDD VSS sg13g2_decap_8
XFILLER_19_770 VDD VSS sg13g2_decap_8
XFILLER_80_334 VDD VSS sg13g2_decap_8
XFILLER_25_217 VDD VSS sg13g2_decap_8
XFILLER_53_559 VDD VSS sg13g2_decap_8
XFILLER_18_280 VDD VSS sg13g2_decap_8
XFILLER_22_924 VDD VSS sg13g2_decap_8
XFILLER_34_784 VDD VSS sg13g2_decap_8
XFILLER_21_434 VDD VSS sg13g2_decap_8
XFILLER_33_294 VDD VSS sg13g2_decap_8
X_1968_ VDD _1968_/Y _1976_/B VSS sg13g2_inv_1
X_1899_ _1899_/B _1899_/A _1903_/A VDD VSS sg13g2_xor2_1
XFILLER_108_35 VDD VSS sg13g2_decap_8
XFILLER_88_401 VDD VSS sg13g2_decap_8
X_2364__284 VDD VSS _2364_/RESET_B sg13g2_tiehi
XFILLER_89_957 VDD VSS sg13g2_decap_4
XFILLER_68_28 VDD VSS sg13g2_decap_8
XFILLER_89_979 VDD VSS sg13g2_fill_1
XFILLER_69_670 VDD VSS sg13g2_decap_4
XFILLER_88_478 VDD VSS sg13g2_decap_8
XFILLER_48_309 VDD VSS sg13g2_fill_2
XFILLER_112_1022 VDD VSS sg13g2_decap_8
XFILLER_69_692 VDD VSS sg13g2_decap_8
XFILLER_57_843 VDD VSS sg13g2_decap_8
XFILLER_57_832 VDD VSS sg13g2_fill_2
XFILLER_84_662 VDD VSS sg13g2_decap_8
XFILLER_84_49 VDD VSS sg13g2_decap_8
XFILLER_57_887 VDD VSS sg13g2_decap_8
XFILLER_29_567 VDD VSS sg13g2_decap_8
XFILLER_17_21 VDD VSS sg13g2_decap_8
XFILLER_17_707 VDD VSS sg13g2_decap_8
XFILLER_44_515 VDD VSS sg13g2_decap_8
XFILLER_72_835 VDD VSS sg13g2_decap_8
XFILLER_83_161 VDD VSS sg13g2_decap_8
XFILLER_16_217 VDD VSS sg13g2_decap_8
XFILLER_17_98 VDD VSS sg13g2_decap_8
XFILLER_71_378 VDD VSS sg13g2_decap_8
XFILLER_25_784 VDD VSS sg13g2_decap_8
XFILLER_13_924 VDD VSS sg13g2_decap_8
XFILLER_40_732 VDD VSS sg13g2_decap_8
XFILLER_12_434 VDD VSS sg13g2_decap_8
XFILLER_9_917 VDD VSS sg13g2_decap_8
XFILLER_33_42 VDD VSS sg13g2_decap_8
XFILLER_24_294 VDD VSS sg13g2_decap_8
XFILLER_32_1001 VDD VSS sg13g2_decap_8
XFILLER_8_427 VDD VSS sg13g2_decap_8
XFILLER_4_644 VDD VSS sg13g2_decap_8
XFILLER_3_154 VDD VSS sg13g2_decap_8
XFILLER_106_594 VDD VSS sg13g2_decap_8
XFILLER_79_412 VDD VSS sg13g2_decap_8
XFILLER_67_607 VDD VSS sg13g2_decap_8
XFILLER_95_938 VDD VSS sg13g2_decap_8
XFILLER_94_426 VDD VSS sg13g2_decap_8
XFILLER_79_489 VDD VSS sg13g2_decap_4
XFILLER_48_821 VDD VSS sg13g2_decap_8
XFILLER_0_861 VDD VSS sg13g2_decap_8
XFILLER_58_72 VDD VSS sg13g2_decap_8
XFILLER_66_139 VDD VSS sg13g2_decap_8
XFILLER_47_331 VDD VSS sg13g2_decap_8
XFILLER_75_651 VDD VSS sg13g2_decap_8
XFILLER_35_504 VDD VSS sg13g2_decap_8
XFILLER_74_161 VDD VSS sg13g2_fill_1
XFILLER_63_846 VDD VSS sg13g2_decap_8
XFILLER_62_323 VDD VSS sg13g2_decap_8
XFILLER_90_654 VDD VSS sg13g2_fill_2
XFILLER_31_721 VDD VSS sg13g2_decap_8
XFILLER_16_784 VDD VSS sg13g2_decap_8
XFILLER_50_518 VDD VSS sg13g2_decap_8
XFILLER_15_294 VDD VSS sg13g2_decap_8
XFILLER_30_231 VDD VSS sg13g2_decap_8
X_1822_ _1878_/A _1930_/A _1822_/B VDD VSS sg13g2_nand2_1
XFILLER_90_70 VDD VSS sg13g2_decap_8
XFILLER_31_798 VDD VSS sg13g2_decap_8
X_1753_ _1741_/Y VDD _1753_/Y VSS _1726_/A _2242_/Q sg13g2_o21ai_1
Xhold427 _2304_/Q VDD VSS hold427/X sg13g2_dlygate4sd3_1
X_1684_ _1719_/A _1692_/A _1723_/A VDD VSS sg13g2_xor2_1
Xhold405 _1330_/Y VDD VSS _1331_/A sg13g2_dlygate4sd3_1
XFILLER_8_994 VDD VSS sg13g2_decap_8
Xhold416 _1237_/Y VDD VSS _2361_/D sg13g2_dlygate4sd3_1
Xhold438 _1651_/Y VDD VSS _1652_/B sg13g2_dlygate4sd3_1
Xhold449 _2210_/Q VDD VSS hold449/X sg13g2_dlygate4sd3_1
XFILLER_48_1030 VDD VSS sg13g2_decap_8
XFILLER_112_553 VDD VSS sg13g2_decap_8
XFILLER_97_242 VDD VSS sg13g2_decap_8
X_2244__255 VDD VSS _2244_/RESET_B sg13g2_tiehi
XFILLER_31_0 VDD VSS sg13g2_decap_8
X_2305_ _2305__91/L_HI VSS VDD _2305_/D _2305_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_85_426 VDD VSS sg13g2_decap_4
XFILLER_85_404 VDD VSS sg13g2_decap_8
X_2236_ _2236_/RESET_B VSS VDD _2236_/D _2236_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_39_843 VDD VSS sg13g2_decap_8
XFILLER_38_320 VDD VSS sg13g2_decap_8
XFILLER_65_150 VDD VSS sg13g2_fill_1
XFILLER_26_504 VDD VSS sg13g2_decap_8
X_2167_ _2167_/RESET_B VSS VDD _2167_/D _2167_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_93_492 VDD VSS sg13g2_fill_1
XFILLER_53_323 VDD VSS sg13g2_decap_4
XFILLER_38_397 VDD VSS sg13g2_decap_8
XFILLER_81_665 VDD VSS sg13g2_decap_4
XFILLER_81_643 VDD VSS sg13g2_fill_1
XFILLER_54_857 VDD VSS sg13g2_decap_8
XFILLER_0_1043 VDD VSS sg13g2_decap_8
X_2098_ _2352_/Q _2351_/Q _2102_/C VDD VSS sg13g2_and2_1
XFILLER_81_687 VDD VSS sg13g2_decap_8
XFILLER_110_14 VDD VSS sg13g2_decap_8
XFILLER_80_164 VDD VSS sg13g2_decap_8
XFILLER_53_389 VDD VSS sg13g2_decap_8
XFILLER_55_1045 VDD VSS sg13g2_decap_8
XFILLER_34_581 VDD VSS sg13g2_decap_8
XFILLER_22_721 VDD VSS sg13g2_decap_8
X_2251__248 VDD VSS _2251_/RESET_B sg13g2_tiehi
XFILLER_16_1029 VDD VSS sg13g2_decap_8
XFILLER_21_231 VDD VSS sg13g2_decap_8
XFILLER_22_798 VDD VSS sg13g2_decap_8
XFILLER_10_938 VDD VSS sg13g2_decap_8
XFILLER_108_815 VDD VSS sg13g2_decap_8
X_2230__80 VDD VSS _2230__80/L_HI sg13g2_tiehi
XFILLER_79_49 VDD VSS sg13g2_decap_8
XFILLER_89_754 VDD VSS sg13g2_decap_4
XFILLER_77_905 VDD VSS sg13g2_decap_8
XFILLER_88_220 VDD VSS sg13g2_fill_1
XFILLER_1_658 VDD VSS sg13g2_decap_8
XFILLER_77_938 VDD VSS sg13g2_decap_4
XFILLER_76_415 VDD VSS sg13g2_decap_8
XFILLER_49_629 VDD VSS sg13g2_decap_8
XFILLER_0_168 VDD VSS sg13g2_decap_8
XFILLER_88_297 VDD VSS sg13g2_decap_8
XFILLER_76_448 VDD VSS sg13g2_decap_8
XFILLER_48_139 VDD VSS sg13g2_decap_8
XFILLER_85_971 VDD VSS sg13g2_decap_4
XFILLER_17_504 VDD VSS sg13g2_decap_8
XFILLER_28_42 VDD VSS sg13g2_decap_8
XFILLER_29_364 VDD VSS sg13g2_decap_8
XFILLER_57_695 VDD VSS sg13g2_decap_8
XFILLER_44_301 VDD VSS sg13g2_decap_8
XFILLER_56_194 VDD VSS sg13g2_decap_8
XFILLER_60_827 VDD VSS sg13g2_decap_8
XFILLER_32_518 VDD VSS sg13g2_decap_8
XFILLER_44_378 VDD VSS sg13g2_decap_8
XFILLER_25_581 VDD VSS sg13g2_decap_8
XFILLER_13_721 VDD VSS sg13g2_decap_8
XFILLER_44_63 VDD VSS sg13g2_decap_8
XFILLER_12_231 VDD VSS sg13g2_decap_8
XFILLER_9_714 VDD VSS sg13g2_decap_8
XFILLER_100_91 VDD VSS sg13g2_decap_8
XFILLER_8_224 VDD VSS sg13g2_decap_8
XFILLER_13_798 VDD VSS sg13g2_decap_8
XFILLER_60_73 VDD VSS sg13g2_decap_8
XFILLER_5_931 VDD VSS sg13g2_decap_8
XFILLER_4_441 VDD VSS sg13g2_decap_8
XFILLER_5_35 VDD VSS sg13g2_decap_8
XFILLER_107_870 VDD VSS sg13g2_decap_8
XFILLER_67_415 VDD VSS sg13g2_decap_8
XFILLER_94_223 VDD VSS sg13g2_fill_1
X_2021_ _1889_/A _1878_/B _2021_/S _2021_/X VDD VSS sg13g2_mux2_1
XFILLER_85_70 VDD VSS sg13g2_decap_8
XFILLER_94_289 VDD VSS sg13g2_decap_8
XFILLER_82_429 VDD VSS sg13g2_decap_8
XFILLER_63_621 VDD VSS sg13g2_decap_8
XFILLER_48_673 VDD VSS sg13g2_decap_8
XFILLER_35_301 VDD VSS sg13g2_decap_8
XFILLER_78_1056 VDD VSS sg13g2_decap_4
XFILLER_39_1018 VDD VSS sg13g2_decap_8
XFILLER_36_868 VDD VSS sg13g2_decap_8
XFILLER_91_985 VDD VSS sg13g2_fill_1
XFILLER_90_462 VDD VSS sg13g2_decap_8
XFILLER_23_518 VDD VSS sg13g2_decap_8
XFILLER_35_378 VDD VSS sg13g2_decap_8
X_2354__272 VDD VSS _2354_/RESET_B sg13g2_tiehi
XFILLER_50_304 VDD VSS sg13g2_decap_8
XFILLER_16_581 VDD VSS sg13g2_decap_8
XFILLER_31_595 VDD VSS sg13g2_decap_8
X_1805_ _1804_/Y VDD _1809_/B VSS _1812_/A _1800_/Y sg13g2_o21ai_1
XFILLER_79_0 VDD VSS sg13g2_decap_8
X_1736_ VSS VDD _1898_/A _1898_/B _1915_/A _1729_/Y sg13g2_a21oi_1
XFILLER_8_791 VDD VSS sg13g2_decap_8
X_1667_ _1670_/A _1667_/B _2305_/D VDD VSS sg13g2_nor2_1
XFILLER_104_328 VDD VSS sg13g2_decap_8
X_1598_ _1633_/A _1606_/A _1637_/A VDD VSS sg13g2_xor2_1
XFILLER_112_350 VDD VSS sg13g2_decap_8
XFILLER_105_14 VDD VSS sg13g2_decap_8
XFILLER_100_545 VDD VSS sg13g2_decap_4
XFILLER_98_595 VDD VSS sg13g2_decap_8
XFILLER_86_746 VDD VSS sg13g2_decap_8
XFILLER_74_919 VDD VSS sg13g2_decap_8
XFILLER_100_567 VDD VSS sg13g2_decap_8
XFILLER_85_245 VDD VSS sg13g2_decap_8
XFILLER_73_407 VDD VSS sg13g2_decap_8
XFILLER_67_971 VDD VSS sg13g2_decap_8
XFILLER_22_1022 VDD VSS sg13g2_decap_8
XFILLER_39_640 VDD VSS sg13g2_decap_8
X_2219_ _2219_/RESET_B VSS VDD _2219_/D _2219_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_66_470 VDD VSS sg13g2_fill_2
XFILLER_38_161 VDD VSS sg13g2_decap_8
XFILLER_26_301 VDD VSS sg13g2_decap_8
XFILLER_82_963 VDD VSS sg13g2_decap_8
XFILLER_81_440 VDD VSS sg13g2_decap_8
XFILLER_54_654 VDD VSS sg13g2_decap_8
XFILLER_54_632 VDD VSS sg13g2_fill_2
XFILLER_42_805 VDD VSS sg13g2_decap_8
XFILLER_27_868 VDD VSS sg13g2_decap_8
XFILLER_54_698 VDD VSS sg13g2_decap_8
XFILLER_14_518 VDD VSS sg13g2_decap_8
XFILLER_26_378 VDD VSS sg13g2_decap_8
XFILLER_41_315 VDD VSS sg13g2_decap_8
XFILLER_81_28 VDD VSS sg13g2_decap_8
XFILLER_22_595 VDD VSS sg13g2_decap_8
XFILLER_14_77 VDD VSS sg13g2_decap_8
XFILLER_10_735 VDD VSS sg13g2_decap_8
XFILLER_108_612 VDD VSS sg13g2_decap_8
XFILLER_6_728 VDD VSS sg13g2_decap_8
XFILLER_30_21 VDD VSS sg13g2_decap_8
XFILLER_107_133 VDD VSS sg13g2_decap_8
XFILLER_5_238 VDD VSS sg13g2_decap_8
XFILLER_108_689 VDD VSS sg13g2_decap_8
XFILLER_30_98 VDD VSS sg13g2_decap_8
XFILLER_2_945 VDD VSS sg13g2_decap_8
XFILLER_89_551 VDD VSS sg13g2_decap_8
XFILLER_77_702 VDD VSS sg13g2_decap_8
XFILLER_1_455 VDD VSS sg13g2_decap_8
Xclk_pad IOVDD IOVSS clk_pad/p2c clk_PAD VDD VSS sg13g2_IOPadIn
XFILLER_77_746 VDD VSS sg13g2_decap_8
XFILLER_103_383 VDD VSS sg13g2_decap_8
XFILLER_76_212 VDD VSS sg13g2_decap_8
XFILLER_39_63 VDD VSS sg13g2_decap_8
XFILLER_49_426 VDD VSS sg13g2_decap_8
XFILLER_92_749 VDD VSS sg13g2_decap_8
XFILLER_76_289 VDD VSS sg13g2_decap_8
XFILLER_17_301 VDD VSS sg13g2_decap_8
XFILLER_29_161 VDD VSS sg13g2_decap_8
XFILLER_73_952 VDD VSS sg13g2_decap_8
XFILLER_91_248 VDD VSS sg13g2_decap_8
XFILLER_18_868 VDD VSS sg13g2_decap_8
XFILLER_44_120 VDD VSS sg13g2_decap_8
XFILLER_73_974 VDD VSS sg13g2_fill_2
XFILLER_72_462 VDD VSS sg13g2_decap_8
XFILLER_33_805 VDD VSS sg13g2_decap_8
XFILLER_17_378 VDD VSS sg13g2_decap_8
XFILLER_55_95 VDD VSS sg13g2_decap_8
XFILLER_32_315 VDD VSS sg13g2_decap_8
XFILLER_44_186 VDD VSS sg13g2_decap_8
XFILLER_41_860 VDD VSS sg13g2_decap_8
XFILLER_9_511 VDD VSS sg13g2_decap_8
XFILLER_13_595 VDD VSS sg13g2_decap_8
XFILLER_40_370 VDD VSS sg13g2_decap_8
XFILLER_72_7 VDD VSS sg13g2_decap_8
XFILLER_9_588 VDD VSS sg13g2_decap_8
XFILLER_99_304 VDD VSS sg13g2_decap_8
X_1521_ _1602_/B _1521_/B _2283_/D VDD VSS sg13g2_and2_1
XFILLER_84_1060 VDD VSS sg13g2_fill_1
X_1452_ VSS VDD _1370_/Y _1453_/B _2245_/D _1451_/Y sg13g2_a21oi_1
XFILLER_101_309 VDD VSS sg13g2_decap_8
X_1383_ _1383_/Y _1383_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_68_757 VDD VSS sg13g2_decap_8
XFILLER_67_223 VDD VSS sg13g2_decap_8
XFILLER_110_865 VDD VSS sg13g2_decap_8
XFILLER_83_705 VDD VSS sg13g2_decap_8
XFILLER_96_91 VDD VSS sg13g2_decap_8
XFILLER_56_919 VDD VSS sg13g2_fill_1
XFILLER_76_790 VDD VSS sg13g2_decap_8
XFILLER_82_215 VDD VSS sg13g2_decap_8
X_2004_ _2071_/B _2004_/B _2004_/Y VDD VSS sg13g2_nor2_1
XFILLER_63_440 VDD VSS sg13g2_decap_8
XFILLER_36_665 VDD VSS sg13g2_decap_8
XFILLER_24_805 VDD VSS sg13g2_decap_8
XFILLER_90_270 VDD VSS sg13g2_decap_8
XFILLER_23_315 VDD VSS sg13g2_decap_8
XFILLER_35_175 VDD VSS sg13g2_decap_8
XFILLER_91_1042 VDD VSS sg13g2_decap_8
XFILLER_52_1004 VDD VSS sg13g2_decap_8
XFILLER_51_668 VDD VSS sg13g2_decap_8
XFILLER_50_134 VDD VSS sg13g2_fill_2
XFILLER_32_882 VDD VSS sg13g2_decap_8
XFILLER_52_1059 VDD VSS sg13g2_fill_2
XFILLER_31_392 VDD VSS sg13g2_decap_8
X_1719_ _1720_/B _1719_/A _1719_/B VDD VSS sg13g2_xnor2_1
XFILLER_105_637 VDD VSS sg13g2_decap_8
XFILLER_104_147 VDD VSS sg13g2_decap_8
XFILLER_101_821 VDD VSS sg13g2_decap_8
XFILLER_76_28 VDD VSS sg13g2_decap_8
XFILLER_59_735 VDD VSS sg13g2_decap_8
XFILLER_58_201 VDD VSS sg13g2_decap_8
XFILLER_101_865 VDD VSS sg13g2_decap_4
XFILLER_101_876 VDD VSS sg13g2_decap_8
XFILLER_74_716 VDD VSS sg13g2_decap_8
XFILLER_47_908 VDD VSS sg13g2_decap_8
XFILLER_58_234 VDD VSS sg13g2_decap_8
XFILLER_46_407 VDD VSS sg13g2_decap_8
XFILLER_86_598 VDD VSS sg13g2_decap_4
XFILLER_100_386 VDD VSS sg13g2_decap_4
XFILLER_73_215 VDD VSS sg13g2_decap_8
XFILLER_39_492 VDD VSS sg13g2_decap_8
XFILLER_82_771 VDD VSS sg13g2_decap_8
XFILLER_92_49 VDD VSS sg13g2_decap_8
XFILLER_55_996 VDD VSS sg13g2_fill_1
XFILLER_42_602 VDD VSS sg13g2_decap_8
XFILLER_27_665 VDD VSS sg13g2_decap_8
XFILLER_15_805 VDD VSS sg13g2_decap_8
XFILLER_25_21 VDD VSS sg13g2_decap_8
XFILLER_70_955 VDD VSS sg13g2_decap_8
XFILLER_81_270 VDD VSS sg13g2_decap_8
XFILLER_54_495 VDD VSS sg13g2_decap_8
XFILLER_14_315 VDD VSS sg13g2_decap_8
XFILLER_41_112 VDD VSS sg13g2_decap_8
XFILLER_26_175 VDD VSS sg13g2_decap_8
XFILLER_42_679 VDD VSS sg13g2_decap_8
XFILLER_30_819 VDD VSS sg13g2_decap_8
XFILLER_23_882 VDD VSS sg13g2_decap_8
XFILLER_25_98 VDD VSS sg13g2_decap_8
XFILLER_109_910 VDD VSS sg13g2_decap_8
XFILLER_10_532 VDD VSS sg13g2_decap_8
XFILLER_22_392 VDD VSS sg13g2_decap_8
XFILLER_6_525 VDD VSS sg13g2_decap_8
XFILLER_41_42 VDD VSS sg13g2_decap_8
XFILLER_109_987 VDD VSS sg13g2_decap_8
XFILLER_108_464 VDD VSS sg13g2_decap_8
X_2264__225 VDD VSS _2264_/RESET_B sg13g2_tiehi
XFILLER_9_0 VDD VSS sg13g2_decap_8
XFILLER_2_742 VDD VSS sg13g2_decap_8
XFILLER_1_252 VDD VSS sg13g2_decap_8
XFILLER_96_329 VDD VSS sg13g2_decap_8
XFILLER_2_14 VDD VSS sg13g2_decap_8
XFILLER_49_212 VDD VSS sg13g2_decap_8
XFILLER_77_565 VDD VSS sg13g2_decap_8
XFILLER_38_919 VDD VSS sg13g2_decap_8
XFILLER_49_267 VDD VSS sg13g2_decap_8
XFILLER_64_226 VDD VSS sg13g2_decap_8
XFILLER_92_579 VDD VSS sg13g2_decap_8
XFILLER_73_782 VDD VSS sg13g2_decap_8
XFILLER_46_996 VDD VSS sg13g2_decap_8
XFILLER_61_900 VDD VSS sg13g2_decap_8
XFILLER_33_602 VDD VSS sg13g2_decap_8
XFILLER_18_665 VDD VSS sg13g2_decap_8
XFILLER_45_462 VDD VSS sg13g2_decap_8
XFILLER_61_944 VDD VSS sg13g2_decap_8
XFILLER_17_175 VDD VSS sg13g2_decap_8
XFILLER_32_112 VDD VSS sg13g2_decap_8
XFILLER_75_1059 VDD VSS sg13g2_fill_2
XFILLER_33_679 VDD VSS sg13g2_decap_8
XFILLER_21_819 VDD VSS sg13g2_decap_8
XFILLER_20_329 VDD VSS sg13g2_decap_8
XFILLER_14_882 VDD VSS sg13g2_decap_8
XFILLER_32_189 VDD VSS sg13g2_decap_8
XFILLER_13_392 VDD VSS sg13g2_decap_8
XFILLER_9_385 VDD VSS sg13g2_decap_8
XFILLER_12_1043 VDD VSS sg13g2_decap_8
XFILLER_99_112 VDD VSS sg13g2_decap_8
X_1504_ _2150_/A VDD _1504_/Y VSS _2110_/A _1503_/X sg13g2_o21ai_1
XFILLER_82_1019 VDD VSS sg13g2_decap_8
XFILLER_99_156 VDD VSS sg13g2_decap_8
X_1435_ VDD _2237_/D _1435_/A VSS sg13g2_inv_1
XFILLER_68_565 VDD VSS sg13g2_decap_8
X_1366_ _2266_/Q _1495_/C _1366_/A _1366_/Y VDD VSS sg13g2_nand3_1
XFILLER_110_662 VDD VSS sg13g2_decap_8
XFILLER_96_885 VDD VSS sg13g2_decap_8
XFILLER_83_502 VDD VSS sg13g2_fill_1
XFILLER_56_749 VDD VSS sg13g2_decap_8
XFILLER_83_557 VDD VSS sg13g2_decap_8
X_1297_ VDD _2178_/D _1297_/A VSS sg13g2_inv_1
XFILLER_37_952 VDD VSS sg13g2_decap_8
XFILLER_49_790 VDD VSS sg13g2_decap_8
XFILLER_64_760 VDD VSS sg13g2_decap_8
XFILLER_24_602 VDD VSS sg13g2_decap_8
XFILLER_55_259 VDD VSS sg13g2_decap_8
XFILLER_36_462 VDD VSS sg13g2_decap_8
XFILLER_70_229 VDD VSS sg13g2_decap_8
XFILLER_52_922 VDD VSS sg13g2_decap_8
XFILLER_23_112 VDD VSS sg13g2_decap_8
XFILLER_24_679 VDD VSS sg13g2_decap_8
XFILLER_51_443 VDD VSS sg13g2_decap_8
XFILLER_12_819 VDD VSS sg13g2_decap_8
XFILLER_51_476 VDD VSS sg13g2_decap_8
XFILLER_11_329 VDD VSS sg13g2_decap_8
XFILLER_23_189 VDD VSS sg13g2_decap_8
XFILLER_108_1060 VDD VSS sg13g2_fill_1
XFILLER_20_896 VDD VSS sg13g2_decap_8
XFILLER_106_902 VDD VSS sg13g2_decap_8
XFILLER_11_56 VDD VSS sg13g2_decap_8
XFILLER_3_539 VDD VSS sg13g2_decap_8
XFILLER_106_979 VDD VSS sg13g2_decap_8
XFILLER_105_456 VDD VSS sg13g2_decap_8
XFILLER_87_49 VDD VSS sg13g2_decap_8
XFILLER_2_7 VDD VSS sg13g2_decap_8
XFILLER_28_1050 VDD VSS sg13g2_decap_8
XFILLER_47_705 VDD VSS sg13g2_decap_8
XFILLER_59_532 VDD VSS sg13g2_decap_8
XFILLER_87_896 VDD VSS sg13g2_decap_8
XFILLER_87_885 VDD VSS sg13g2_decap_8
XFILLER_86_384 VDD VSS sg13g2_decap_8
XFILLER_4_1008 VDD VSS sg13g2_decap_8
XFILLER_28_952 VDD VSS sg13g2_decap_8
XFILLER_62_719 VDD VSS sg13g2_decap_8
XFILLER_15_602 VDD VSS sg13g2_decap_8
XFILLER_36_42 VDD VSS sg13g2_decap_8
XFILLER_27_462 VDD VSS sg13g2_decap_8
XFILLER_82_590 VDD VSS sg13g2_decap_8
XFILLER_43_933 VDD VSS sg13g2_decap_8
XFILLER_14_112 VDD VSS sg13g2_decap_8
XFILLER_70_752 VDD VSS sg13g2_decap_8
XFILLER_54_292 VDD VSS sg13g2_decap_8
XFILLER_15_679 VDD VSS sg13g2_decap_8
XFILLER_42_454 VDD VSS sg13g2_decap_8
XFILLER_30_616 VDD VSS sg13g2_decap_8
XFILLER_14_189 VDD VSS sg13g2_decap_8
XFILLER_35_1043 VDD VSS sg13g2_decap_8
XFILLER_7_812 VDD VSS sg13g2_decap_8
XFILLER_52_96 VDD VSS sg13g2_decap_4
XFILLER_6_322 VDD VSS sg13g2_decap_8
XFILLER_11_896 VDD VSS sg13g2_decap_8
XFILLER_109_784 VDD VSS sg13g2_decap_8
XFILLER_108_250 VDD VSS sg13g2_decap_8
XFILLER_7_889 VDD VSS sg13g2_decap_8
XFILLER_6_399 VDD VSS sg13g2_decap_8
XFILLER_112_938 VDD VSS sg13g2_decap_8
XFILLER_81_1041 VDD VSS sg13g2_decap_8
XFILLER_96_126 VDD VSS sg13g2_decap_8
XFILLER_35_7 VDD VSS sg13g2_decap_8
XFILLER_78_874 VDD VSS sg13g2_decap_8
XFILLER_78_841 VDD VSS sg13g2_decap_4
XFILLER_111_448 VDD VSS sg13g2_decap_8
X_1220_ _1220_/A _2352_/Q _2099_/B _1221_/B VDD VSS sg13g2_nor3_1
XFILLER_93_811 VDD VSS sg13g2_decap_8
XFILLER_77_384 VDD VSS sg13g2_decap_8
XFILLER_42_1036 VDD VSS sg13g2_decap_8
XFILLER_38_716 VDD VSS sg13g2_decap_8
XFILLER_93_866 VDD VSS sg13g2_decap_8
XFILLER_65_557 VDD VSS sg13g2_decap_8
XFILLER_19_952 VDD VSS sg13g2_decap_8
XFILLER_92_354 VDD VSS sg13g2_decap_8
XFILLER_80_516 VDD VSS sg13g2_decap_8
XFILLER_18_462 VDD VSS sg13g2_decap_8
XFILLER_37_259 VDD VSS sg13g2_decap_8
XFILLER_93_70 VDD VSS sg13g2_decap_8
XFILLER_46_782 VDD VSS sg13g2_decap_8
XFILLER_34_966 VDD VSS sg13g2_decap_8
XFILLER_21_616 VDD VSS sg13g2_decap_8
XFILLER_33_476 VDD VSS sg13g2_decap_8
X_1984_ _1988_/A _1984_/A _1984_/B VDD VSS sg13g2_xnor2_1
XFILLER_60_284 VDD VSS sg13g2_decap_8
XFILLER_20_126 VDD VSS sg13g2_decap_8
XFILLER_9_182 VDD VSS sg13g2_decap_8
XFILLER_61_0 VDD VSS sg13g2_decap_8
XFILLER_103_938 VDD VSS sg13g2_decap_8
XFILLER_88_649 VDD VSS sg13g2_fill_2
XFILLER_69_830 VDD VSS sg13g2_decap_8
X_1418_ _1418_/Y _1418_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_87_137 VDD VSS sg13g2_decap_8
XFILLER_68_340 VDD VSS sg13g2_decap_8
XFILLER_96_693 VDD VSS sg13g2_decap_8
X_1349_ VDD _2203_/D _1349_/A VSS sg13g2_inv_1
XFILLER_56_546 VDD VSS sg13g2_fill_1
XFILLER_29_749 VDD VSS sg13g2_decap_8
XFILLER_84_899 VDD VSS sg13g2_decap_8
XFILLER_71_516 VDD VSS sg13g2_fill_2
XFILLER_28_259 VDD VSS sg13g2_decap_8
XFILLER_25_966 VDD VSS sg13g2_decap_8
XFILLER_40_914 VDD VSS sg13g2_decap_8
XFILLER_12_616 VDD VSS sg13g2_decap_8
XFILLER_24_476 VDD VSS sg13g2_decap_8
XFILLER_51_251 VDD VSS sg13g2_decap_8
XFILLER_11_126 VDD VSS sg13g2_decap_8
XFILLER_8_609 VDD VSS sg13g2_decap_8
X_2330__189 VDD VSS _2330_/RESET_B sg13g2_tiehi
XFILLER_7_119 VDD VSS sg13g2_decap_8
XIO_BOND_vss_pads\[0\].vss_pad VSS bondpad_70x70
XFILLER_20_693 VDD VSS sg13g2_decap_8
XFILLER_4_826 VDD VSS sg13g2_decap_8
XFILLER_22_77 VDD VSS sg13g2_decap_8
XFILLER_3_336 VDD VSS sg13g2_decap_8
XFILLER_106_776 VDD VSS sg13g2_decap_8
XFILLER_105_242 VDD VSS sg13g2_decap_8
XFILLER_65_1036 VDD VSS sg13g2_decap_8
XFILLER_79_638 VDD VSS sg13g2_decap_8
XFILLER_78_126 VDD VSS sg13g2_decap_8
XFILLER_94_608 VDD VSS sg13g2_decap_8
XFILLER_87_682 VDD VSS sg13g2_decap_8
XFILLER_59_362 VDD VSS sg13g2_decap_8
XFILLER_47_502 VDD VSS sg13g2_decap_8
XFILLER_75_855 VDD VSS sg13g2_decap_8
XFILLER_86_192 VDD VSS sg13g2_decap_8
XFILLER_74_321 VDD VSS sg13g2_decap_8
XFILLER_47_63 VDD VSS sg13g2_decap_8
XFILLER_47_557 VDD VSS sg13g2_decap_8
XFILLER_19_259 VDD VSS sg13g2_decap_8
XFILLER_90_858 VDD VSS sg13g2_decap_8
XFILLER_103_91 VDD VSS sg13g2_decap_8
XFILLER_43_730 VDD VSS sg13g2_decap_8
XFILLER_31_903 VDD VSS sg13g2_decap_8
XFILLER_16_966 VDD VSS sg13g2_decap_8
XFILLER_72_1018 VDD VSS sg13g2_decap_8
XFILLER_15_476 VDD VSS sg13g2_decap_8
XFILLER_30_413 VDD VSS sg13g2_decap_8
XFILLER_42_273 VDD VSS sg13g2_decap_8
XFILLER_8_35 VDD VSS sg13g2_decap_8
XFILLER_11_693 VDD VSS sg13g2_decap_8
XFILLER_109_581 VDD VSS sg13g2_decap_8
XFILLER_7_686 VDD VSS sg13g2_decap_8
XFILLER_6_196 VDD VSS sg13g2_decap_8
XFILLER_112_735 VDD VSS sg13g2_decap_8
X_2321_ _2321_/RESET_B VSS VDD _2321_/D _2321_/Q _2337_/CLK sg13g2_dfrbpq_1
XFILLER_88_70 VDD VSS sg13g2_decap_8
XFILLER_111_245 VDD VSS sg13g2_decap_8
XFILLER_69_148 VDD VSS sg13g2_fill_2
X_2252_ _2252_/RESET_B VSS VDD _2252_/D _2252_/Q clkload0/A sg13g2_dfrbpq_1
X_2203__134 VDD VSS _2203_/RESET_B sg13g2_tiehi
X_1203_ VDD _1222_/B _2093_/A VSS sg13g2_inv_1
XFILLER_38_502 VDD VSS sg13g2_decap_8
X_2183_ _2183_/RESET_B VSS VDD _2183_/D _2183_/Q _2371_/CLK sg13g2_dfrbpq_1
XFILLER_53_505 VDD VSS sg13g2_decap_8
XFILLER_80_313 VDD VSS sg13g2_decap_8
XFILLER_53_516 VDD VSS sg13g2_fill_1
XFILLER_22_903 VDD VSS sg13g2_decap_8
XFILLER_34_763 VDD VSS sg13g2_decap_8
XFILLER_21_413 VDD VSS sg13g2_decap_8
XFILLER_33_273 VDD VSS sg13g2_decap_8
X_1967_ _1967_/B _1967_/A _1976_/B VDD VSS sg13g2_xor2_1
XFILLER_30_980 VDD VSS sg13g2_decap_8
XFILLER_88_1047 VDD VSS sg13g2_decap_8
XFILLER_88_1014 VDD VSS sg13g2_decap_4
XFILLER_107_507 VDD VSS sg13g2_decap_8
X_1898_ _1898_/B _1898_/A _1899_/B VDD VSS sg13g2_xor2_1
XFILLER_108_14 VDD VSS sg13g2_decap_8
XFILLER_89_936 VDD VSS sg13g2_decap_8
XFILLER_102_223 VDD VSS sg13g2_fill_2
XFILLER_102_234 VDD VSS sg13g2_decap_8
XFILLER_88_457 VDD VSS sg13g2_decap_8
XFILLER_57_800 VDD VSS sg13g2_decap_8
XFILLER_112_1001 VDD VSS sg13g2_decap_8
XFILLER_97_991 VDD VSS sg13g2_decap_8
XFILLER_84_641 VDD VSS sg13g2_decap_8
XFILLER_84_28 VDD VSS sg13g2_decap_8
XFILLER_29_546 VDD VSS sg13g2_decap_8
XFILLER_72_814 VDD VSS sg13g2_decap_8
XFILLER_56_354 VDD VSS sg13g2_decap_4
XFILLER_95_1029 VDD VSS sg13g2_decap_8
XFILLER_56_398 VDD VSS sg13g2_decap_8
XFILLER_71_357 VDD VSS sg13g2_decap_8
XFILLER_17_77 VDD VSS sg13g2_decap_8
XFILLER_40_711 VDD VSS sg13g2_decap_8
XFILLER_25_763 VDD VSS sg13g2_decap_8
XFILLER_13_903 VDD VSS sg13g2_decap_8
XFILLER_12_413 VDD VSS sg13g2_decap_8
XFILLER_33_21 VDD VSS sg13g2_decap_8
XFILLER_24_273 VDD VSS sg13g2_decap_8
XFILLER_71_1040 VDD VSS sg13g2_decap_8
XFILLER_40_788 VDD VSS sg13g2_decap_8
XFILLER_8_406 VDD VSS sg13g2_decap_8
XFILLER_21_980 VDD VSS sg13g2_decap_8
XFILLER_33_98 VDD VSS sg13g2_decap_8
XFILLER_32_1057 VDD VSS sg13g2_decap_4
XFILLER_20_490 VDD VSS sg13g2_decap_8
XFILLER_4_623 VDD VSS sg13g2_decap_8
XFILLER_109_0 VDD VSS sg13g2_decap_8
XFILLER_3_133 VDD VSS sg13g2_decap_8
XFILLER_106_573 VDD VSS sg13g2_decap_8
XFILLER_95_917 VDD VSS sg13g2_decap_8
XFILLER_0_840 VDD VSS sg13g2_decap_8
XFILLER_94_405 VDD VSS sg13g2_decap_8
XFILLER_79_468 VDD VSS sg13g2_decap_8
XFILLER_48_800 VDD VSS sg13g2_decap_8
XFILLER_75_630 VDD VSS sg13g2_decap_8
XFILLER_74_140 VDD VSS sg13g2_decap_8
XFILLER_48_877 VDD VSS sg13g2_decap_8
XFILLER_90_622 VDD VSS sg13g2_decap_8
XFILLER_63_825 VDD VSS sg13g2_decap_8
XFILLER_62_302 VDD VSS sg13g2_decap_8
XFILLER_31_700 VDD VSS sg13g2_decap_8
XFILLER_62_379 VDD VSS sg13g2_decap_8
XFILLER_16_763 VDD VSS sg13g2_decap_8
XFILLER_15_273 VDD VSS sg13g2_decap_8
XFILLER_30_210 VDD VSS sg13g2_decap_8
X_1821_ VSS VDD _1822_/B _1821_/B _1889_/A sg13g2_or2_1
XFILLER_31_777 VDD VSS sg13g2_decap_8
XFILLER_12_980 VDD VSS sg13g2_decap_8
XFILLER_30_287 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_10_clk clkbuf_leaf_9_clk/A _2337_/CLK VDD VSS sg13g2_buf_8
X_1752_ VSS VDD _1761_/A _1751_/B _1752_/Y _1749_/A sg13g2_a21oi_1
XFILLER_11_490 VDD VSS sg13g2_decap_8
XFILLER_8_973 VDD VSS sg13g2_decap_8
X_1683_ _1719_/A _2319_/Q _2305_/Q VDD VSS sg13g2_xnor2_1
Xhold406 _2260_/Q VDD VSS _2110_/B sg13g2_dlygate4sd3_1
Xhold417 _2209_/Q VDD VSS hold417/X sg13g2_dlygate4sd3_1
XFILLER_7_483 VDD VSS sg13g2_decap_8
Xhold428 _1663_/Y VDD VSS _1664_/B sg13g2_dlygate4sd3_1
XFILLER_99_91 VDD VSS sg13g2_decap_8
Xhold439 _2289_/Q VDD VSS _1594_/A sg13g2_dlygate4sd3_1
XFILLER_98_711 VDD VSS sg13g2_decap_8
XFILLER_112_532 VDD VSS sg13g2_decap_8
XFILLER_97_221 VDD VSS sg13g2_decap_8
X_2304_ _2304__95/L_HI VSS VDD _2304_/D _2304_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_98_799 VDD VSS sg13g2_decap_8
XFILLER_24_0 VDD VSS sg13g2_decap_8
XFILLER_100_738 VDD VSS sg13g2_fill_2
X_2235_ _2235_/RESET_B VSS VDD _2235_/D _2235_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_66_630 VDD VSS sg13g2_decap_8
XFILLER_39_822 VDD VSS sg13g2_decap_8
XFILLER_57_129 VDD VSS sg13g2_decap_8
X_2166_ _2166_/RESET_B VSS VDD _2166_/D _2166_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_94_983 VDD VSS sg13g2_decap_8
XFILLER_81_622 VDD VSS sg13g2_decap_8
XFILLER_54_836 VDD VSS sg13g2_decap_8
XFILLER_39_899 VDD VSS sg13g2_decap_8
XFILLER_38_376 VDD VSS sg13g2_decap_8
XFILLER_80_143 VDD VSS sg13g2_decap_8
XFILLER_65_184 VDD VSS sg13g2_decap_8
XFILLER_0_1022 VDD VSS sg13g2_decap_8
X_2097_ VSS VDD _2099_/B _2095_/Y _2351_/D _2096_/Y sg13g2_a21oi_1
XFILLER_34_560 VDD VSS sg13g2_decap_8
XFILLER_22_700 VDD VSS sg13g2_decap_8
XFILLER_53_368 VDD VSS sg13g2_decap_8
XFILLER_0_91 VDD VSS sg13g2_decap_8
XFILLER_55_1024 VDD VSS sg13g2_decap_8
XFILLER_61_390 VDD VSS sg13g2_decap_8
XFILLER_16_1008 VDD VSS sg13g2_decap_8
XFILLER_21_210 VDD VSS sg13g2_decap_8
XFILLER_22_777 VDD VSS sg13g2_decap_8
XFILLER_10_917 VDD VSS sg13g2_decap_8
XFILLER_21_287 VDD VSS sg13g2_decap_8
XFILLER_102_7 VDD VSS sg13g2_decap_8
XFILLER_79_28 VDD VSS sg13g2_decap_8
XFILLER_103_510 VDD VSS sg13g2_decap_8
XFILLER_62_1006 VDD VSS sg13g2_decap_4
XFILLER_1_637 VDD VSS sg13g2_decap_8
XFILLER_88_276 VDD VSS sg13g2_decap_8
XFILLER_0_147 VDD VSS sg13g2_decap_8
XFILLER_95_49 VDD VSS sg13g2_decap_8
XFILLER_28_21 VDD VSS sg13g2_decap_8
XFILLER_48_118 VDD VSS sg13g2_decap_8
XFILLER_85_950 VDD VSS sg13g2_decap_8
XFILLER_29_343 VDD VSS sg13g2_decap_8
XFILLER_72_622 VDD VSS sg13g2_fill_1
XFILLER_57_674 VDD VSS sg13g2_decap_8
XFILLER_56_173 VDD VSS sg13g2_decap_8
XFILLER_28_98 VDD VSS sg13g2_decap_8
XFILLER_72_655 VDD VSS sg13g2_decap_8
XFILLER_60_806 VDD VSS sg13g2_decap_8
XFILLER_45_869 VDD VSS sg13g2_decap_8
XFILLER_44_357 VDD VSS sg13g2_decap_8
XFILLER_71_176 VDD VSS sg13g2_decap_8
XFILLER_25_560 VDD VSS sg13g2_decap_8
XFILLER_13_700 VDD VSS sg13g2_decap_8
XFILLER_44_42 VDD VSS sg13g2_decap_8
XFILLER_71_198 VDD VSS sg13g2_decap_8
XFILLER_53_880 VDD VSS sg13g2_decap_8
XFILLER_12_210 VDD VSS sg13g2_decap_8
XFILLER_8_203 VDD VSS sg13g2_decap_8
XFILLER_13_777 VDD VSS sg13g2_decap_8
XFILLER_100_70 VDD VSS sg13g2_decap_8
XFILLER_40_585 VDD VSS sg13g2_decap_8
XFILLER_12_287 VDD VSS sg13g2_decap_8
XFILLER_60_52 VDD VSS sg13g2_decap_8
XFILLER_5_910 VDD VSS sg13g2_decap_8
XFILLER_4_420 VDD VSS sg13g2_decap_8
XFILLER_5_14 VDD VSS sg13g2_decap_8
XFILLER_5_987 VDD VSS sg13g2_decap_8
XFILLER_79_232 VDD VSS sg13g2_fill_2
XFILLER_79_210 VDD VSS sg13g2_decap_8
XFILLER_4_497 VDD VSS sg13g2_decap_8
XFILLER_95_714 VDD VSS sg13g2_decap_8
XFILLER_79_243 VDD VSS sg13g2_decap_8
X_2020_ _2025_/A _2019_/X _2020_/Y VDD VSS sg13g2_nor2b_1
XFILLER_94_268 VDD VSS sg13g2_decap_4
XFILLER_82_408 VDD VSS sg13g2_decap_8
XFILLER_48_652 VDD VSS sg13g2_decap_8
X_2274__205 VDD VSS _2274_/RESET_B sg13g2_tiehi
XFILLER_78_1035 VDD VSS sg13g2_decap_8
XFILLER_75_493 VDD VSS sg13g2_fill_2
XFILLER_36_847 VDD VSS sg13g2_decap_8
XFILLER_47_184 VDD VSS sg13g2_decap_8
XFILLER_63_677 VDD VSS sg13g2_decap_8
XFILLER_51_839 VDD VSS sg13g2_fill_1
XFILLER_51_828 VDD VSS sg13g2_decap_8
XFILLER_16_560 VDD VSS sg13g2_decap_8
XFILLER_35_357 VDD VSS sg13g2_decap_8
XFILLER_62_176 VDD VSS sg13g2_decap_4
XFILLER_31_574 VDD VSS sg13g2_decap_8
X_1804_ VSS VDD _1800_/C _1802_/Y _1804_/Y _1803_/Y sg13g2_a21oi_1
XFILLER_102_1055 VDD VSS sg13g2_decap_4
X_1735_ _1898_/B _2229_/Q _2237_/Q VDD VSS sg13g2_xnor2_1
XFILLER_8_770 VDD VSS sg13g2_decap_8
XFILLER_105_819 VDD VSS sg13g2_decap_8
XFILLER_7_280 VDD VSS sg13g2_decap_8
X_1666_ _1666_/Y _1646_/Y _1665_/X hold424/X _1189_/Y VDD VSS sg13g2_a22oi_1
XFILLER_104_307 VDD VSS sg13g2_decap_8
X_1597_ _1633_/A _2296_/Q _2281_/Q VDD VSS sg13g2_xnor2_1
XFILLER_98_574 VDD VSS sg13g2_decap_8
XFILLER_100_524 VDD VSS sg13g2_decap_8
XFILLER_85_224 VDD VSS sg13g2_decap_8
XFILLER_67_950 VDD VSS sg13g2_decap_8
XFILLER_22_1001 VDD VSS sg13g2_decap_8
X_2218_ _2218_/RESET_B VSS VDD _2218_/D _2218_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_696 VDD VSS sg13g2_decap_8
XFILLER_38_140 VDD VSS sg13g2_decap_8
XFILLER_82_942 VDD VSS sg13g2_decap_8
X_2149_ _2149_/A _2149_/B _2375_/D VDD VSS sg13g2_and2_1
XFILLER_27_847 VDD VSS sg13g2_decap_8
XFILLER_26_357 VDD VSS sg13g2_decap_8
XFILLER_81_496 VDD VSS sg13g2_decap_8
XFILLER_50_850 VDD VSS sg13g2_decap_8
XFILLER_50_894 VDD VSS sg13g2_fill_1
XFILLER_22_574 VDD VSS sg13g2_decap_8
XFILLER_14_56 VDD VSS sg13g2_decap_8
XFILLER_10_714 VDD VSS sg13g2_decap_8
XFILLER_6_707 VDD VSS sg13g2_decap_8
XFILLER_107_112 VDD VSS sg13g2_decap_8
XFILLER_5_217 VDD VSS sg13g2_decap_8
XFILLER_108_668 VDD VSS sg13g2_decap_8
XFILLER_2_924 VDD VSS sg13g2_decap_8
XFILLER_30_77 VDD VSS sg13g2_decap_8
XFILLER_89_530 VDD VSS sg13g2_decap_8
XFILLER_1_434 VDD VSS sg13g2_decap_8
XFILLER_39_42 VDD VSS sg13g2_decap_8
XFILLER_49_405 VDD VSS sg13g2_decap_8
XFILLER_103_362 VDD VSS sg13g2_decap_8
XFILLER_76_268 VDD VSS sg13g2_decap_8
XFILLER_58_950 VDD VSS sg13g2_decap_4
XFILLER_65_909 VDD VSS sg13g2_decap_8
XFILLER_92_728 VDD VSS sg13g2_decap_8
XFILLER_91_227 VDD VSS sg13g2_decap_8
XFILLER_58_994 VDD VSS sg13g2_decap_8
XFILLER_57_460 VDD VSS sg13g2_decap_4
XFILLER_29_140 VDD VSS sg13g2_decap_8
XFILLER_85_791 VDD VSS sg13g2_decap_8
XFILLER_57_493 VDD VSS sg13g2_decap_8
XFILLER_18_847 VDD VSS sg13g2_decap_8
XFILLER_17_357 VDD VSS sg13g2_decap_8
XFILLER_55_63 VDD VSS sg13g2_decap_8
XFILLER_111_91 VDD VSS sg13g2_decap_8
XFILLER_38_1052 VDD VSS sg13g2_decap_8
XFILLER_71_73 VDD VSS sg13g2_decap_8
XFILLER_13_574 VDD VSS sg13g2_decap_8
XFILLER_9_567 VDD VSS sg13g2_decap_8
XFILLER_65_7 VDD VSS sg13g2_decap_8
XFILLER_5_784 VDD VSS sg13g2_decap_8
X_1520_ _1589_/A hold522/X _1521_/B VDD VSS sg13g2_nor2b_1
X_1451_ _1451_/A _1453_/B _1451_/Y VDD VSS sg13g2_nor2_1
XFILLER_4_294 VDD VSS sg13g2_decap_8
X_1382_ _1382_/Y _1382_/A _1465_/C VDD VSS sg13g2_nand2_1
XFILLER_110_844 VDD VSS sg13g2_decap_8
XFILLER_95_522 VDD VSS sg13g2_decap_8
XFILLER_96_70 VDD VSS sg13g2_decap_8
XFILLER_45_1045 VDD VSS sg13g2_decap_8
XFILLER_67_202 VDD VSS sg13g2_decap_8
XFILLER_95_555 VDD VSS sg13g2_fill_2
X_2003_ _2005_/D _2003_/A _2003_/B VDD VSS sg13g2_xnor2_1
XFILLER_36_644 VDD VSS sg13g2_decap_8
XFILLER_64_986 VDD VSS sg13g2_decap_8
XFILLER_35_154 VDD VSS sg13g2_decap_8
XFILLER_91_794 VDD VSS sg13g2_decap_8
XFILLER_51_647 VDD VSS sg13g2_decap_8
XFILLER_63_496 VDD VSS sg13g2_decap_4
XFILLER_50_113 VDD VSS sg13g2_decap_8
XFILLER_91_1021 VDD VSS sg13g2_decap_8
XFILLER_91_0 VDD VSS sg13g2_decap_8
XFILLER_32_861 VDD VSS sg13g2_decap_8
XFILLER_31_371 VDD VSS sg13g2_decap_8
X_1718_ _1725_/A _1718_/B _1718_/Y VDD VSS sg13g2_nor2_1
XFILLER_105_616 VDD VSS sg13g2_decap_8
XFILLER_104_126 VDD VSS sg13g2_decap_8
X_1649_ _1671_/C _1649_/B _2299_/D VDD VSS sg13g2_nor2_1
XFILLER_101_800 VDD VSS sg13g2_decap_8
XFILLER_99_850 VDD VSS sg13g2_decap_8
XFILLER_98_360 VDD VSS sg13g2_decap_8
XFILLER_58_224 VDD VSS sg13g2_fill_1
XFILLER_101_844 VDD VSS sg13g2_fill_1
XFILLER_100_321 VDD VSS sg13g2_decap_8
XFILLER_86_577 VDD VSS sg13g2_decap_8
XFILLER_55_920 VDD VSS sg13g2_fill_2
XFILLER_6_1050 VDD VSS sg13g2_decap_8
XFILLER_39_471 VDD VSS sg13g2_decap_8
XFILLER_27_644 VDD VSS sg13g2_decap_8
XFILLER_92_28 VDD VSS sg13g2_decap_8
XFILLER_26_154 VDD VSS sg13g2_decap_8
XFILLER_70_934 VDD VSS sg13g2_decap_8
XFILLER_54_474 VDD VSS sg13g2_decap_8
XFILLER_42_658 VDD VSS sg13g2_decap_8
XFILLER_23_861 VDD VSS sg13g2_decap_8
XFILLER_25_77 VDD VSS sg13g2_decap_8
XFILLER_10_511 VDD VSS sg13g2_decap_8
XFILLER_22_371 VDD VSS sg13g2_decap_8
XFILLER_41_21 VDD VSS sg13g2_decap_8
XFILLER_6_504 VDD VSS sg13g2_decap_8
XFILLER_109_966 VDD VSS sg13g2_decap_8
XFILLER_108_443 VDD VSS sg13g2_decap_8
XFILLER_10_588 VDD VSS sg13g2_decap_8
XFILLER_41_98 VDD VSS sg13g2_decap_8
XFILLER_29_1029 VDD VSS sg13g2_decap_8
XFILLER_2_721 VDD VSS sg13g2_decap_8
XFILLER_96_308 VDD VSS sg13g2_decap_8
XFILLER_1_231 VDD VSS sg13g2_decap_8
XFILLER_104_682 VDD VSS sg13g2_decap_8
XFILLER_2_798 VDD VSS sg13g2_decap_8
XFILLER_77_544 VDD VSS sg13g2_decap_8
XFILLER_49_246 VDD VSS sg13g2_decap_8
XFILLER_106_91 VDD VSS sg13g2_decap_8
XFILLER_65_717 VDD VSS sg13g2_decap_8
XFILLER_64_205 VDD VSS sg13g2_decap_8
XFILLER_92_558 VDD VSS sg13g2_decap_8
XFILLER_57_290 VDD VSS sg13g2_decap_8
XFILLER_18_644 VDD VSS sg13g2_decap_8
XFILLER_66_84 VDD VSS sg13g2_decap_8
XFILLER_46_975 VDD VSS sg13g2_decap_8
XFILLER_17_154 VDD VSS sg13g2_decap_8
XFILLER_33_658 VDD VSS sg13g2_decap_8
XFILLER_60_477 VDD VSS sg13g2_decap_8
XFILLER_60_488 VDD VSS sg13g2_fill_2
XFILLER_20_308 VDD VSS sg13g2_decap_8
XFILLER_14_861 VDD VSS sg13g2_decap_8
XFILLER_32_168 VDD VSS sg13g2_decap_8
XFILLER_13_371 VDD VSS sg13g2_decap_8
XFILLER_9_364 VDD VSS sg13g2_decap_8
XFILLER_12_1022 VDD VSS sg13g2_decap_8
X_1503_ _1514_/A _1518_/B _1518_/C _1518_/D _1503_/X VDD VSS sg13g2_and4_1
XFILLER_5_581 VDD VSS sg13g2_decap_8
XFILLER_88_809 VDD VSS sg13g2_decap_8
X_1434_ _1435_/A _1429_/Y hold447/X _1429_/B _1373_/A VDD VSS sg13g2_a22oi_1
XFILLER_110_641 VDD VSS sg13g2_decap_8
XFILLER_96_864 VDD VSS sg13g2_decap_8
XFILLER_68_544 VDD VSS sg13g2_decap_8
X_1365_ _1495_/C _2265_/Q _1365_/B _2355_/Q VDD VSS sg13g2_and3_1
XFILLER_95_385 VDD VSS sg13g2_decap_8
XFILLER_56_728 VDD VSS sg13g2_decap_8
X_1296_ _1296_/Y _1344_/B1 hold332/X _1344_/A2 _2342_/Q VDD VSS sg13g2_a22oi_1
XFILLER_83_536 VDD VSS sg13g2_decap_8
XFILLER_37_931 VDD VSS sg13g2_decap_8
XFILLER_55_238 VDD VSS sg13g2_decap_8
XFILLER_52_901 VDD VSS sg13g2_decap_8
XFILLER_36_441 VDD VSS sg13g2_decap_8
XFILLER_91_591 VDD VSS sg13g2_decap_8
XFILLER_102_49 VDD VSS sg13g2_decap_8
XFILLER_51_422 VDD VSS sg13g2_decap_8
XFILLER_24_658 VDD VSS sg13g2_decap_8
X_2213__114 VDD VSS _2213_/RESET_B sg13g2_tiehi
XFILLER_11_308 VDD VSS sg13g2_decap_8
XFILLER_23_168 VDD VSS sg13g2_decap_8
XFILLER_20_875 VDD VSS sg13g2_decap_8
XFILLER_3_518 VDD VSS sg13g2_decap_8
XFILLER_11_35 VDD VSS sg13g2_decap_8
XFILLER_106_958 VDD VSS sg13g2_decap_8
XFILLER_105_435 VDD VSS sg13g2_decap_8
XFILLER_87_28 VDD VSS sg13g2_decap_8
XFILLER_99_680 VDD VSS sg13g2_decap_8
XFILLER_59_511 VDD VSS sg13g2_decap_8
XFILLER_87_864 VDD VSS sg13g2_decap_8
XFILLER_98_190 VDD VSS sg13g2_decap_8
XFILLER_101_685 VDD VSS sg13g2_decap_8
XFILLER_86_363 VDD VSS sg13g2_decap_8
XFILLER_74_514 VDD VSS sg13g2_fill_1
XFILLER_100_140 VDD VSS sg13g2_decap_8
XFILLER_100_173 VDD VSS sg13g2_fill_2
XFILLER_100_184 VDD VSS sg13g2_decap_8
XFILLER_74_525 VDD VSS sg13g2_fill_2
XFILLER_28_931 VDD VSS sg13g2_decap_8
XFILLER_36_21 VDD VSS sg13g2_decap_8
XFILLER_46_227 VDD VSS sg13g2_decap_8
XFILLER_43_912 VDD VSS sg13g2_decap_8
XFILLER_27_441 VDD VSS sg13g2_decap_8
XFILLER_70_731 VDD VSS sg13g2_decap_8
XFILLER_55_783 VDD VSS sg13g2_decap_8
XFILLER_15_658 VDD VSS sg13g2_decap_8
XFILLER_36_98 VDD VSS sg13g2_decap_8
XFILLER_42_433 VDD VSS sg13g2_decap_8
XFILLER_43_989 VDD VSS sg13g2_decap_8
XFILLER_35_1022 VDD VSS sg13g2_decap_8
XFILLER_14_168 VDD VSS sg13g2_decap_8
XFILLER_52_75 VDD VSS sg13g2_decap_8
XFILLER_6_301 VDD VSS sg13g2_decap_8
XFILLER_11_875 VDD VSS sg13g2_decap_8
XFILLER_10_385 VDD VSS sg13g2_decap_8
XFILLER_7_868 VDD VSS sg13g2_decap_8
XFILLER_109_763 VDD VSS sg13g2_decap_8
XFILLER_6_378 VDD VSS sg13g2_decap_8
XFILLER_112_917 VDD VSS sg13g2_decap_8
XFILLER_105_980 VDD VSS sg13g2_decap_8
XFILLER_78_820 VDD VSS sg13g2_decap_8
XFILLER_111_427 VDD VSS sg13g2_decap_8
XFILLER_96_105 VDD VSS sg13g2_decap_8
XFILLER_42_1015 VDD VSS sg13g2_decap_8
XFILLER_2_595 VDD VSS sg13g2_decap_8
XFILLER_28_7 VDD VSS sg13g2_decap_8
XFILLER_92_333 VDD VSS sg13g2_decap_8
XFILLER_65_536 VDD VSS sg13g2_decap_8
XFILLER_19_931 VDD VSS sg13g2_decap_8
XFILLER_37_238 VDD VSS sg13g2_decap_8
XFILLER_46_761 VDD VSS sg13g2_decap_8
XFILLER_18_441 VDD VSS sg13g2_decap_8
XFILLER_34_945 VDD VSS sg13g2_decap_8
XFILLER_33_455 VDD VSS sg13g2_decap_8
XFILLER_60_263 VDD VSS sg13g2_decap_8
XFILLER_20_105 VDD VSS sg13g2_decap_8
X_1983_ _1995_/A _1995_/B _2000_/C VDD VSS sg13g2_nor2_1
XFILLER_9_161 VDD VSS sg13g2_decap_8
XFILLER_54_0 VDD VSS sg13g2_decap_8
XFILLER_103_917 VDD VSS sg13g2_decap_8
XFILLER_88_628 VDD VSS sg13g2_decap_8
XFILLER_87_116 VDD VSS sg13g2_decap_8
XFILLER_102_449 VDD VSS sg13g2_decap_8
X_1417_ _1416_/Y VDD _2229_/D VSS _1373_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_96_672 VDD VSS sg13g2_decap_8
XFILLER_69_875 VDD VSS sg13g2_fill_2
XFILLER_29_728 VDD VSS sg13g2_decap_8
XFILLER_68_363 VDD VSS sg13g2_fill_1
XFILLER_3_91 VDD VSS sg13g2_decap_8
XFILLER_111_994 VDD VSS sg13g2_decap_8
XFILLER_95_182 VDD VSS sg13g2_decap_8
X_1348_ _1349_/A _1347_/Y hold537/X _1347_/B _1364_/A VDD VSS sg13g2_a22oi_1
XFILLER_28_238 VDD VSS sg13g2_decap_8
X_1279_ VDD _2169_/D _1279_/A VSS sg13g2_inv_1
XFILLER_84_878 VDD VSS sg13g2_decap_8
XFILLER_25_945 VDD VSS sg13g2_decap_8
XFILLER_51_230 VDD VSS sg13g2_decap_8
Xin_data_pads\[2\].in_data_pad IOVDD IOVSS _1373_/A in_data_PADs[2] VDD VSS sg13g2_IOPadIn
XFILLER_11_105 VDD VSS sg13g2_decap_8
XFILLER_24_455 VDD VSS sg13g2_decap_8
XFILLER_20_672 VDD VSS sg13g2_decap_8
XFILLER_22_56 VDD VSS sg13g2_decap_8
XFILLER_4_805 VDD VSS sg13g2_decap_8
XFILLER_98_49 VDD VSS sg13g2_decap_8
XFILLER_3_315 VDD VSS sg13g2_decap_8
XFILLER_106_755 VDD VSS sg13g2_decap_8
XFILLER_105_221 VDD VSS sg13g2_decap_8
XFILLER_65_1015 VDD VSS sg13g2_decap_8
XFILLER_79_617 VDD VSS sg13g2_decap_8
XFILLER_78_105 VDD VSS sg13g2_decap_8
X_2261__229 VDD VSS _2261_/RESET_B sg13g2_tiehi
XFILLER_93_119 VDD VSS sg13g2_decap_8
XFILLER_59_341 VDD VSS sg13g2_decap_8
XFILLER_75_834 VDD VSS sg13g2_decap_8
XFILLER_86_171 VDD VSS sg13g2_decap_8
XFILLER_74_300 VDD VSS sg13g2_decap_8
XFILLER_19_238 VDD VSS sg13g2_decap_8
XFILLER_47_42 VDD VSS sg13g2_decap_8
XFILLER_74_366 VDD VSS sg13g2_decap_8
XFILLER_103_70 VDD VSS sg13g2_decap_8
XFILLER_16_945 VDD VSS sg13g2_decap_8
XFILLER_43_786 VDD VSS sg13g2_decap_8
XFILLER_15_455 VDD VSS sg13g2_decap_8
XFILLER_63_63 VDD VSS sg13g2_decap_8
XFILLER_42_252 VDD VSS sg13g2_decap_8
XFILLER_31_959 VDD VSS sg13g2_decap_8
XFILLER_8_14 VDD VSS sg13g2_decap_8
XFILLER_30_469 VDD VSS sg13g2_decap_8
XFILLER_11_672 VDD VSS sg13g2_decap_8
XFILLER_109_560 VDD VSS sg13g2_decap_8
XFILLER_10_182 VDD VSS sg13g2_decap_8
XFILLER_7_665 VDD VSS sg13g2_decap_8
XFILLER_6_175 VDD VSS sg13g2_decap_8
XFILLER_112_714 VDD VSS sg13g2_decap_8
XFILLER_97_414 VDD VSS sg13g2_decap_8
X_2320_ _2320_/RESET_B VSS VDD _2320_/D _2320_/Q clkload9/A sg13g2_dfrbpq_1
XFILLER_3_882 VDD VSS sg13g2_decap_8
XFILLER_111_224 VDD VSS sg13g2_decap_8
XFILLER_69_127 VDD VSS sg13g2_decap_8
X_2251_ _2251_/RESET_B VSS VDD _2251_/D _2251_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_2_392 VDD VSS sg13g2_decap_8
XFILLER_84_119 VDD VSS sg13g2_decap_8
X_1202_ VDD _2106_/A _1236_/C VSS sg13g2_inv_1
X_2182_ _2182_/RESET_B VSS VDD _2182_/D _2182_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_78_683 VDD VSS sg13g2_decap_8
XFILLER_77_182 VDD VSS sg13g2_decap_8
XFILLER_93_642 VDD VSS sg13g2_decap_8
XFILLER_81_815 VDD VSS sg13g2_decap_4
XFILLER_38_569 VDD VSS sg13g2_decap_8
XFILLER_92_185 VDD VSS sg13g2_decap_8
XFILLER_65_399 VDD VSS sg13g2_decap_8
XFILLER_34_742 VDD VSS sg13g2_decap_8
XFILLER_80_369 VDD VSS sg13g2_decap_8
XFILLER_61_561 VDD VSS sg13g2_fill_1
XFILLER_61_550 VDD VSS sg13g2_decap_8
XFILLER_33_252 VDD VSS sg13g2_decap_8
XFILLER_22_959 VDD VSS sg13g2_decap_8
XFILLER_61_583 VDD VSS sg13g2_decap_8
X_1966_ _1966_/A _1966_/B _1976_/A VDD VSS sg13g2_nor2_1
XFILLER_18_1050 VDD VSS sg13g2_decap_8
XFILLER_21_469 VDD VSS sg13g2_decap_8
X_1897_ VDD _1973_/A _1897_/A VSS sg13g2_inv_1
XFILLER_89_915 VDD VSS sg13g2_decap_8
XFILLER_1_819 VDD VSS sg13g2_decap_8
XFILLER_88_436 VDD VSS sg13g2_decap_8
XFILLER_0_329 VDD VSS sg13g2_decap_8
XFILLER_25_1043 VDD VSS sg13g2_decap_8
XFILLER_111_791 VDD VSS sg13g2_decap_8
XFILLER_84_620 VDD VSS sg13g2_decap_8
XFILLER_75_119 VDD VSS sg13g2_decap_8
XFILLER_29_525 VDD VSS sg13g2_decap_8
XFILLER_112_1057 VDD VSS sg13g2_decap_4
XFILLER_56_333 VDD VSS sg13g2_decap_8
XFILLER_95_1008 VDD VSS sg13g2_decap_8
XFILLER_84_697 VDD VSS sg13g2_fill_2
XFILLER_56_377 VDD VSS sg13g2_decap_8
XFILLER_17_56 VDD VSS sg13g2_decap_8
XFILLER_83_185 VDD VSS sg13g2_decap_8
XFILLER_25_742 VDD VSS sg13g2_decap_8
XFILLER_80_870 VDD VSS sg13g2_fill_1
XFILLER_24_252 VDD VSS sg13g2_decap_8
XFILLER_52_583 VDD VSS sg13g2_decap_8
XFILLER_13_959 VDD VSS sg13g2_decap_8
XFILLER_40_767 VDD VSS sg13g2_decap_8
XFILLER_12_469 VDD VSS sg13g2_decap_8
XFILLER_33_77 VDD VSS sg13g2_decap_8
XFILLER_32_1036 VDD VSS sg13g2_decap_8
XFILLER_4_602 VDD VSS sg13g2_decap_8
XFILLER_3_112 VDD VSS sg13g2_decap_8
XFILLER_4_679 VDD VSS sg13g2_decap_8
XFILLER_79_447 VDD VSS sg13g2_decap_8
XFILLER_3_189 VDD VSS sg13g2_decap_8
XFILLER_102_780 VDD VSS sg13g2_decap_8
XFILLER_0_896 VDD VSS sg13g2_decap_8
XFILLER_66_119 VDD VSS sg13g2_decap_8
XFILLER_101_290 VDD VSS sg13g2_decap_8
XFILLER_63_804 VDD VSS sg13g2_decap_8
XFILLER_90_601 VDD VSS sg13g2_decap_8
XFILLER_75_686 VDD VSS sg13g2_decap_8
XFILLER_35_539 VDD VSS sg13g2_decap_8
XFILLER_74_84 VDD VSS sg13g2_decap_8
XFILLER_62_358 VDD VSS sg13g2_fill_1
XFILLER_16_742 VDD VSS sg13g2_decap_8
XFILLER_47_399 VDD VSS sg13g2_decap_8
XFILLER_90_689 VDD VSS sg13g2_decap_8
XFILLER_15_252 VDD VSS sg13g2_decap_8
XFILLER_71_881 VDD VSS sg13g2_fill_2
XFILLER_95_7 VDD VSS sg13g2_decap_8
XFILLER_43_583 VDD VSS sg13g2_decap_8
X_1820_ _1889_/B _1930_/A _1821_/B VDD VSS sg13g2_nand2_1
XFILLER_31_756 VDD VSS sg13g2_decap_8
XFILLER_30_266 VDD VSS sg13g2_decap_8
X_1751_ _1761_/A _1751_/B _1751_/X VDD VSS sg13g2_and2_1
XFILLER_8_952 VDD VSS sg13g2_decap_8
Xhold407 _2254_/Q VDD VSS _1199_/A sg13g2_dlygate4sd3_1
X_1682_ _1692_/A _2320_/Q _2306_/Q VDD VSS sg13g2_xnor2_1
Xhold418 _1360_/Y VDD VSS _1361_/A sg13g2_dlygate4sd3_1
XFILLER_7_462 VDD VSS sg13g2_decap_8
XFILLER_99_70 VDD VSS sg13g2_decap_8
Xhold429 _2299_/Q VDD VSS _1685_/B sg13g2_dlygate4sd3_1
XFILLER_112_511 VDD VSS sg13g2_decap_8
XFILLER_97_200 VDD VSS sg13g2_decap_8
X_2303_ _2303__99/L_HI VSS VDD _2303_/D _2303_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_100_717 VDD VSS sg13g2_decap_8
XFILLER_98_778 VDD VSS sg13g2_decap_8
XFILLER_97_277 VDD VSS sg13g2_decap_8
XFILLER_58_609 VDD VSS sg13g2_decap_8
XFILLER_39_801 VDD VSS sg13g2_decap_8
XFILLER_57_108 VDD VSS sg13g2_decap_8
XFILLER_112_588 VDD VSS sg13g2_decap_8
XFILLER_97_288 VDD VSS sg13g2_fill_2
X_2234_ _2234_/RESET_B VSS VDD _2234_/D _2234_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_94_962 VDD VSS sg13g2_decap_8
X_2165_ _2165_/RESET_B VSS VDD _2165_/D _2165_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_39_878 VDD VSS sg13g2_decap_8
XFILLER_17_0 VDD VSS sg13g2_decap_8
XFILLER_65_141 VDD VSS sg13g2_decap_8
XFILLER_38_355 VDD VSS sg13g2_decap_8
XFILLER_81_601 VDD VSS sg13g2_decap_8
XFILLER_93_483 VDD VSS sg13g2_decap_8
XFILLER_54_815 VDD VSS sg13g2_decap_8
XFILLER_0_1001 VDD VSS sg13g2_decap_8
XFILLER_65_163 VDD VSS sg13g2_decap_8
XFILLER_0_70 VDD VSS sg13g2_decap_8
XFILLER_26_539 VDD VSS sg13g2_decap_8
X_2096_ _2107_/B1 VDD _2096_/Y VSS _2099_/B _2102_/B sg13g2_o21ai_1
XFILLER_94_1041 VDD VSS sg13g2_decap_8
XFILLER_41_509 VDD VSS sg13g2_decap_8
XFILLER_80_199 VDD VSS sg13g2_decap_8
XFILLER_110_49 VDD VSS sg13g2_decap_8
XFILLER_62_892 VDD VSS sg13g2_decap_8
XFILLER_22_756 VDD VSS sg13g2_decap_8
XFILLER_21_266 VDD VSS sg13g2_decap_8
X_1949_ _1949_/B _1949_/A _1951_/B VDD VSS sg13g2_xor2_1
XFILLER_107_305 VDD VSS sg13g2_decap_8
XFILLER_1_616 VDD VSS sg13g2_decap_8
XFILLER_103_544 VDD VSS sg13g2_decap_8
XFILLER_0_126 VDD VSS sg13g2_decap_8
XFILLER_88_255 VDD VSS sg13g2_decap_8
XFILLER_95_28 VDD VSS sg13g2_decap_8
XFILLER_103_588 VDD VSS sg13g2_decap_8
XFILLER_69_480 VDD VSS sg13g2_decap_8
XFILLER_57_653 VDD VSS sg13g2_decap_8
XFILLER_29_322 VDD VSS sg13g2_decap_8
XFILLER_28_77 VDD VSS sg13g2_decap_8
XFILLER_56_152 VDD VSS sg13g2_decap_8
XFILLER_72_634 VDD VSS sg13g2_decap_8
XFILLER_71_111 VDD VSS sg13g2_decap_8
XFILLER_17_539 VDD VSS sg13g2_decap_8
XFILLER_29_399 VDD VSS sg13g2_decap_8
XFILLER_44_336 VDD VSS sg13g2_decap_8
XFILLER_72_689 VDD VSS sg13g2_fill_1
XFILLER_72_667 VDD VSS sg13g2_decap_4
XFILLER_71_155 VDD VSS sg13g2_decap_8
XFILLER_44_21 VDD VSS sg13g2_decap_8
XFILLER_52_391 VDD VSS sg13g2_fill_1
XFILLER_13_756 VDD VSS sg13g2_decap_8
XFILLER_40_564 VDD VSS sg13g2_decap_8
XFILLER_12_266 VDD VSS sg13g2_decap_8
XFILLER_9_749 VDD VSS sg13g2_decap_8
XFILLER_60_31 VDD VSS sg13g2_fill_1
XFILLER_8_259 VDD VSS sg13g2_decap_8
XFILLER_5_966 VDD VSS sg13g2_decap_8
XFILLER_109_91 VDD VSS sg13g2_decap_8
XFILLER_4_476 VDD VSS sg13g2_decap_8
XFILLER_106_393 VDD VSS sg13g2_decap_8
XFILLER_79_266 VDD VSS sg13g2_decap_4
XFILLER_94_203 VDD VSS sg13g2_decap_8
XFILLER_39_119 VDD VSS sg13g2_decap_8
XFILLER_94_247 VDD VSS sg13g2_decap_8
XFILLER_48_631 VDD VSS sg13g2_decap_8
XFILLER_10_7 VDD VSS sg13g2_decap_8
XFILLER_0_693 VDD VSS sg13g2_decap_8
XFILLER_78_1014 VDD VSS sg13g2_decap_8
XFILLER_76_984 VDD VSS sg13g2_decap_8
XFILLER_75_472 VDD VSS sg13g2_decap_8
XFILLER_36_826 VDD VSS sg13g2_decap_8
XFILLER_91_954 VDD VSS sg13g2_fill_2
XFILLER_63_656 VDD VSS sg13g2_decap_8
XFILLER_35_336 VDD VSS sg13g2_decap_8
XFILLER_51_807 VDD VSS sg13g2_decap_8
XFILLER_62_155 VDD VSS sg13g2_decap_8
XFILLER_90_497 VDD VSS sg13g2_decap_8
XFILLER_62_199 VDD VSS sg13g2_decap_8
XFILLER_50_339 VDD VSS sg13g2_decap_8
XFILLER_31_553 VDD VSS sg13g2_decap_8
X_1803_ _1797_/Y VDD _1803_/Y VSS _1776_/A _2226_/Q sg13g2_o21ai_1
XFILLER_102_1034 VDD VSS sg13g2_decap_8
X_1734_ _1730_/Y VDD _1898_/A VSS _1926_/A _1732_/Y sg13g2_o21ai_1
XFILLER_85_1029 VDD VSS sg13g2_decap_8
X_1665_ _2310_/Q _2334_/Q _2326_/Q _2349_/Q _2341_/Q _1677_/A _1665_/X VDD VSS sg13g2_mux4_1
X_1596_ _1606_/A _2297_/Q _2282_/Q VDD VSS sg13g2_xnor2_1
XFILLER_98_553 VDD VSS sg13g2_decap_8
XFILLER_59_929 VDD VSS sg13g2_decap_8
XFILLER_58_406 VDD VSS sg13g2_decap_8
XFILLER_112_385 VDD VSS sg13g2_decap_8
XFILLER_100_503 VDD VSS sg13g2_decap_8
XFILLER_61_1040 VDD VSS sg13g2_decap_8
X_2217_ _2217_/RESET_B VSS VDD _2217_/D _2217_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_105_49 VDD VSS sg13g2_decap_8
XFILLER_82_921 VDD VSS sg13g2_decap_8
XFILLER_22_1057 VDD VSS sg13g2_decap_4
XFILLER_39_675 VDD VSS sg13g2_decap_8
XFILLER_27_826 VDD VSS sg13g2_decap_8
XFILLER_66_472 VDD VSS sg13g2_fill_1
X_2148_ _2149_/A _2148_/B _2374_/D VDD VSS sg13g2_and2_1
XFILLER_53_111 VDD VSS sg13g2_decap_8
XFILLER_53_122 VDD VSS sg13g2_fill_1
XFILLER_26_336 VDD VSS sg13g2_decap_8
XFILLER_38_196 VDD VSS sg13g2_decap_8
XFILLER_82_998 VDD VSS sg13g2_decap_8
X_2079_ _2069_/X _2086_/A _2079_/S _2080_/B VDD VSS sg13g2_mux2_1
XFILLER_81_475 VDD VSS sg13g2_decap_8
XFILLER_50_840 VDD VSS sg13g2_decap_4
XFILLER_22_553 VDD VSS sg13g2_decap_8
XFILLER_14_35 VDD VSS sg13g2_decap_8
XFILLER_50_873 VDD VSS sg13g2_decap_8
XFILLER_108_647 VDD VSS sg13g2_decap_8
XFILLER_30_56 VDD VSS sg13g2_decap_8
XFILLER_107_168 VDD VSS sg13g2_decap_8
XFILLER_2_903 VDD VSS sg13g2_decap_8
XFILLER_104_820 VDD VSS sg13g2_decap_8
XFILLER_1_413 VDD VSS sg13g2_decap_8
XFILLER_103_341 VDD VSS sg13g2_decap_8
XFILLER_39_21 VDD VSS sg13g2_decap_8
XFILLER_76_203 VDD VSS sg13g2_decap_4
XFILLER_7_1029 VDD VSS sg13g2_decap_8
XFILLER_76_247 VDD VSS sg13g2_decap_8
XFILLER_39_98 VDD VSS sg13g2_decap_8
XFILLER_85_770 VDD VSS sg13g2_decap_8
XFILLER_91_206 VDD VSS sg13g2_decap_8
XFILLER_58_973 VDD VSS sg13g2_decap_8
XFILLER_64_409 VDD VSS sg13g2_fill_2
XFILLER_18_826 VDD VSS sg13g2_decap_8
XFILLER_17_336 VDD VSS sg13g2_decap_8
XFILLER_55_42 VDD VSS sg13g2_decap_8
XFILLER_29_196 VDD VSS sg13g2_decap_8
XFILLER_73_998 VDD VSS sg13g2_fill_2
XFILLER_72_497 VDD VSS sg13g2_decap_8
XFILLER_38_1031 VDD VSS sg13g2_decap_8
XFILLER_111_70 VDD VSS sg13g2_decap_8
XFILLER_13_553 VDD VSS sg13g2_decap_8
XFILLER_71_63 VDD VSS sg13g2_fill_1
XFILLER_41_895 VDD VSS sg13g2_decap_8
XFILLER_9_546 VDD VSS sg13g2_decap_8
XFILLER_5_763 VDD VSS sg13g2_decap_8
XFILLER_58_7 VDD VSS sg13g2_decap_8
XFILLER_84_1051 VDD VSS sg13g2_decap_8
XFILLER_99_339 VDD VSS sg13g2_decap_8
X_1450_ VSS VDD _1364_/Y _1455_/B _2244_/D _1449_/Y sg13g2_a21oi_1
XFILLER_4_273 VDD VSS sg13g2_decap_8
X_1381_ _1380_/Y VDD _2215_/D VSS _1367_/B _1379_/Y sg13g2_o21ai_1
XFILLER_45_1024 VDD VSS sg13g2_decap_8
XFILLER_68_715 VDD VSS sg13g2_decap_8
XFILLER_110_823 VDD VSS sg13g2_decap_8
XFILLER_1_980 VDD VSS sg13g2_decap_8
XFILLER_67_258 VDD VSS sg13g2_decap_8
XFILLER_0_490 VDD VSS sg13g2_decap_8
XFILLER_95_589 VDD VSS sg13g2_decap_8
XFILLER_49_995 VDD VSS sg13g2_decap_8
X_2002_ _2025_/A _2071_/A _2089_/S VDD VSS sg13g2_nand2_1
XFILLER_36_623 VDD VSS sg13g2_decap_8
XFILLER_91_773 VDD VSS sg13g2_decap_8
XFILLER_64_976 VDD VSS sg13g2_fill_2
XFILLER_64_965 VDD VSS sg13g2_decap_8
XFILLER_35_133 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_91_1000 VDD VSS sg13g2_decap_8
XFILLER_51_626 VDD VSS sg13g2_decap_8
XFILLER_63_475 VDD VSS sg13g2_decap_8
XFILLER_32_840 VDD VSS sg13g2_decap_8
X_2174__192 VDD VSS _2174_/RESET_B sg13g2_tiehi
XFILLER_50_158 VDD VSS sg13g2_decap_8
XFILLER_31_350 VDD VSS sg13g2_decap_8
XFILLER_84_0 VDD VSS sg13g2_decap_8
X_1717_ _1716_/Y VDD _1717_/Y VSS _1724_/S hold539/X sg13g2_o21ai_1
XFILLER_104_105 VDD VSS sg13g2_decap_8
X_1648_ _1648_/Y _1646_/Y _1647_/X _1685_/B _1671_/B VDD VSS sg13g2_a22oi_1
XFILLER_6_91 VDD VSS sg13g2_decap_8
XFILLER_100_300 VDD VSS sg13g2_decap_8
XFILLER_98_383 VDD VSS sg13g2_decap_8
X_1579_ VSS VDD _1580_/A1 _1207_/Y _1579_/Y _1522_/Y sg13g2_a21oi_1
XFILLER_86_556 VDD VSS sg13g2_decap_8
XFILLER_112_182 VDD VSS sg13g2_decap_8
XFILLER_39_450 VDD VSS sg13g2_decap_8
XFILLER_55_954 VDD VSS sg13g2_fill_1
XFILLER_55_943 VDD VSS sg13g2_decap_8
XFILLER_67_792 VDD VSS sg13g2_fill_1
XFILLER_27_623 VDD VSS sg13g2_decap_8
XFILLER_82_751 VDD VSS sg13g2_decap_8
XFILLER_70_913 VDD VSS sg13g2_decap_8
XFILLER_55_987 VDD VSS sg13g2_decap_8
XFILLER_54_453 VDD VSS sg13g2_decap_8
XFILLER_26_133 VDD VSS sg13g2_decap_8
XFILLER_42_637 VDD VSS sg13g2_decap_8
XFILLER_109_1029 VDD VSS sg13g2_decap_8
XFILLER_23_840 VDD VSS sg13g2_decap_8
XFILLER_25_56 VDD VSS sg13g2_decap_8
X_2333__177 VDD VSS _2333_/RESET_B sg13g2_tiehi
XFILLER_22_350 VDD VSS sg13g2_decap_8
XFILLER_50_692 VDD VSS sg13g2_fill_2
XFILLER_10_567 VDD VSS sg13g2_decap_8
XFILLER_109_945 VDD VSS sg13g2_decap_8
XFILLER_108_422 VDD VSS sg13g2_decap_8
XFILLER_41_77 VDD VSS sg13g2_decap_8
XFILLER_2_700 VDD VSS sg13g2_decap_8
XFILLER_29_1008 VDD VSS sg13g2_decap_8
XFILLER_1_210 VDD VSS sg13g2_decap_8
XFILLER_111_609 VDD VSS sg13g2_decap_8
XFILLER_104_661 VDD VSS sg13g2_decap_8
XFILLER_77_523 VDD VSS sg13g2_decap_8
XFILLER_110_119 VDD VSS sg13g2_decap_8
XFILLER_2_777 VDD VSS sg13g2_decap_8
XFILLER_49_203 VDD VSS sg13g2_decap_4
XFILLER_103_182 VDD VSS sg13g2_decap_8
XFILLER_106_70 VDD VSS sg13g2_decap_8
XFILLER_1_287 VDD VSS sg13g2_decap_8
XFILLER_2_49 VDD VSS sg13g2_decap_8
XFILLER_66_63 VDD VSS sg13g2_decap_8
XFILLER_92_526 VDD VSS sg13g2_decap_8
XFILLER_46_954 VDD VSS sg13g2_decap_8
XFILLER_58_781 VDD VSS sg13g2_decap_8
XFILLER_18_623 VDD VSS sg13g2_decap_8
XFILLER_73_751 VDD VSS sg13g2_fill_1
XFILLER_17_133 VDD VSS sg13g2_decap_8
XFILLER_75_1017 VDD VSS sg13g2_fill_2
XFILLER_72_250 VDD VSS sg13g2_decap_4
XFILLER_33_637 VDD VSS sg13g2_decap_8
XFILLER_60_412 VDD VSS sg13g2_decap_8
XFILLER_45_497 VDD VSS sg13g2_decap_8
XFILLER_72_294 VDD VSS sg13g2_decap_8
XFILLER_82_84 VDD VSS sg13g2_decap_8
XFILLER_60_456 VDD VSS sg13g2_decap_4
XFILLER_14_840 VDD VSS sg13g2_decap_8
XFILLER_32_147 VDD VSS sg13g2_decap_8
XFILLER_13_350 VDD VSS sg13g2_decap_8
XFILLER_41_692 VDD VSS sg13g2_decap_8
XFILLER_9_343 VDD VSS sg13g2_decap_8
XFILLER_12_1001 VDD VSS sg13g2_decap_8
X_1502_ _1502_/A _2093_/A _2150_/B _1502_/D _1518_/D VDD VSS sg13g2_nor4_1
XFILLER_5_560 VDD VSS sg13g2_decap_8
XFILLER_102_609 VDD VSS sg13g2_decap_8
XFILLER_99_147 VDD VSS sg13g2_decap_4
X_1433_ VDD _2236_/D _1433_/A VSS sg13g2_inv_1
XFILLER_101_119 VDD VSS sg13g2_decap_8
XFILLER_68_501 VDD VSS sg13g2_decap_8
XFILLER_110_620 VDD VSS sg13g2_decap_8
XFILLER_96_843 VDD VSS sg13g2_decap_8
XFILLER_95_342 VDD VSS sg13g2_decap_8
X_1364_ _1364_/Y _1364_/A _1465_/C VDD VSS sg13g2_nand2_1
X_1295_ VDD _2177_/D _1295_/A VSS sg13g2_inv_1
XFILLER_56_707 VDD VSS sg13g2_decap_8
XFILLER_37_910 VDD VSS sg13g2_decap_8
XFILLER_110_697 VDD VSS sg13g2_decap_8
XFILLER_55_217 VDD VSS sg13g2_decap_8
XFILLER_36_420 VDD VSS sg13g2_decap_8
XFILLER_102_28 VDD VSS sg13g2_decap_8
XFILLER_37_987 VDD VSS sg13g2_decap_8
XFILLER_91_570 VDD VSS sg13g2_decap_8
XFILLER_64_795 VDD VSS sg13g2_decap_8
XFILLER_24_637 VDD VSS sg13g2_decap_8
XFILLER_36_497 VDD VSS sg13g2_decap_8
XFILLER_63_283 VDD VSS sg13g2_decap_8
XFILLER_23_147 VDD VSS sg13g2_decap_8
XFILLER_20_854 VDD VSS sg13g2_decap_8
XFILLER_11_14 VDD VSS sg13g2_decap_8
XFILLER_106_937 VDD VSS sg13g2_decap_8
XFILLER_105_414 VDD VSS sg13g2_decap_8
XFILLER_78_309 VDD VSS sg13g2_decap_4
XFILLER_87_843 VDD VSS sg13g2_decap_8
XFILLER_86_342 VDD VSS sg13g2_decap_8
XFILLER_59_567 VDD VSS sg13g2_decap_8
XFILLER_28_910 VDD VSS sg13g2_decap_8
XFILLER_46_206 VDD VSS sg13g2_decap_8
XFILLER_98_1039 VDD VSS sg13g2_decap_8
XFILLER_27_420 VDD VSS sg13g2_decap_8
XFILLER_39_280 VDD VSS sg13g2_decap_4
XFILLER_55_762 VDD VSS sg13g2_decap_8
XFILLER_70_710 VDD VSS sg13g2_decap_8
XFILLER_28_987 VDD VSS sg13g2_decap_8
XFILLER_36_77 VDD VSS sg13g2_decap_8
XFILLER_42_412 VDD VSS sg13g2_decap_8
XFILLER_43_968 VDD VSS sg13g2_decap_8
XFILLER_15_637 VDD VSS sg13g2_decap_8
XFILLER_27_497 VDD VSS sg13g2_decap_8
XFILLER_70_787 VDD VSS sg13g2_decap_8
XFILLER_35_1001 VDD VSS sg13g2_decap_8
XFILLER_14_147 VDD VSS sg13g2_decap_8
XFILLER_52_21 VDD VSS sg13g2_fill_2
XFILLER_11_854 VDD VSS sg13g2_decap_8
XFILLER_109_742 VDD VSS sg13g2_decap_8
XFILLER_10_364 VDD VSS sg13g2_decap_8
XFILLER_7_847 VDD VSS sg13g2_decap_8
XFILLER_6_357 VDD VSS sg13g2_decap_8
XFILLER_111_406 VDD VSS sg13g2_decap_8
XFILLER_69_309 VDD VSS sg13g2_decap_8
XFILLER_2_574 VDD VSS sg13g2_decap_8
XFILLER_104_491 VDD VSS sg13g2_decap_8
XFILLER_77_84 VDD VSS sg13g2_decap_8
XFILLER_65_515 VDD VSS sg13g2_decap_8
XFILLER_92_312 VDD VSS sg13g2_decap_8
XFILLER_19_910 VDD VSS sg13g2_decap_8
XFILLER_37_217 VDD VSS sg13g2_decap_8
XFILLER_46_740 VDD VSS sg13g2_decap_8
XFILLER_18_420 VDD VSS sg13g2_decap_8
XFILLER_92_389 VDD VSS sg13g2_decap_8
XFILLER_34_924 VDD VSS sg13g2_decap_8
XFILLER_61_721 VDD VSS sg13g2_decap_8
XFILLER_19_987 VDD VSS sg13g2_decap_8
XFILLER_45_250 VDD VSS sg13g2_decap_4
XFILLER_52_209 VDD VSS sg13g2_decap_8
XFILLER_18_497 VDD VSS sg13g2_decap_8
XFILLER_33_434 VDD VSS sg13g2_decap_8
XFILLER_61_765 VDD VSS sg13g2_decap_8
XFILLER_60_242 VDD VSS sg13g2_decap_8
X_1982_ _1995_/B _1982_/A _1982_/B _1982_/C VDD VSS sg13g2_and3_1
XFILLER_9_140 VDD VSS sg13g2_decap_8
XFILLER_88_607 VDD VSS sg13g2_decap_8
XFILLER_47_0 VDD VSS sg13g2_decap_8
XFILLER_102_428 VDD VSS sg13g2_decap_8
X_1416_ _1416_/Y _1416_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_111_973 VDD VSS sg13g2_decap_8
XFILLER_96_651 VDD VSS sg13g2_decap_8
XFILLER_29_707 VDD VSS sg13g2_decap_8
X_1347_ _2101_/A _1347_/B _1347_/Y VDD VSS sg13g2_nor2_1
XFILLER_56_504 VDD VSS sg13g2_decap_4
XFILLER_3_70 VDD VSS sg13g2_decap_8
XFILLER_110_494 VDD VSS sg13g2_decap_8
XFILLER_95_161 VDD VSS sg13g2_decap_8
XFILLER_56_526 VDD VSS sg13g2_decap_8
XFILLER_28_217 VDD VSS sg13g2_decap_8
X_1278_ _1278_/Y _1280_/B1 hold375/X _1280_/A2 _2319_/Q VDD VSS sg13g2_a22oi_1
XFILLER_3_1043 VDD VSS sg13g2_decap_8
XFILLER_97_1050 VDD VSS sg13g2_decap_8
XFILLER_71_518 VDD VSS sg13g2_fill_1
XFILLER_71_529 VDD VSS sg13g2_decap_8
XFILLER_58_1001 VDD VSS sg13g2_decap_8
XFILLER_25_924 VDD VSS sg13g2_decap_8
XFILLER_37_784 VDD VSS sg13g2_decap_8
XFILLER_64_592 VDD VSS sg13g2_decap_8
XFILLER_24_434 VDD VSS sg13g2_decap_8
XFILLER_36_294 VDD VSS sg13g2_decap_8
XFILLER_52_765 VDD VSS sg13g2_decap_8
XFILLER_19_1029 VDD VSS sg13g2_decap_8
XFILLER_40_949 VDD VSS sg13g2_decap_8
XFILLER_20_651 VDD VSS sg13g2_decap_8
XFILLER_22_35 VDD VSS sg13g2_decap_8
XFILLER_106_734 VDD VSS sg13g2_decap_8
XFILLER_98_28 VDD VSS sg13g2_decap_8
XFILLER_105_277 VDD VSS sg13g2_decap_4
XFILLER_87_651 VDD VSS sg13g2_decap_8
XFILLER_87_662 VDD VSS sg13g2_fill_1
XFILLER_47_21 VDD VSS sg13g2_decap_8
XFILLER_102_984 VDD VSS sg13g2_fill_2
XFILLER_101_472 VDD VSS sg13g2_decap_8
XFILLER_59_397 VDD VSS sg13g2_decap_8
XFILLER_19_217 VDD VSS sg13g2_decap_8
XFILLER_74_345 VDD VSS sg13g2_decap_8
XFILLER_41_1060 VDD VSS sg13g2_fill_1
XFILLER_47_98 VDD VSS sg13g2_decap_4
XFILLER_90_827 VDD VSS sg13g2_decap_4
XFILLER_74_389 VDD VSS sg13g2_decap_8
XFILLER_28_784 VDD VSS sg13g2_decap_8
XFILLER_16_924 VDD VSS sg13g2_decap_8
XFILLER_55_581 VDD VSS sg13g2_decap_8
XFILLER_15_434 VDD VSS sg13g2_decap_8
XFILLER_63_42 VDD VSS sg13g2_decap_8
XFILLER_27_294 VDD VSS sg13g2_decap_8
XFILLER_43_765 VDD VSS sg13g2_decap_8
XFILLER_63_75 VDD VSS sg13g2_decap_4
XFILLER_42_231 VDD VSS sg13g2_decap_8
XFILLER_70_584 VDD VSS sg13g2_decap_8
XFILLER_31_938 VDD VSS sg13g2_decap_8
XFILLER_63_97 VDD VSS sg13g2_decap_8
XFILLER_11_651 VDD VSS sg13g2_decap_8
XFILLER_30_448 VDD VSS sg13g2_decap_8
XFILLER_10_161 VDD VSS sg13g2_decap_8
XFILLER_7_644 VDD VSS sg13g2_decap_8
XFILLER_6_154 VDD VSS sg13g2_decap_8
XFILLER_98_905 VDD VSS sg13g2_fill_2
XFILLER_98_938 VDD VSS sg13g2_decap_8
XFILLER_111_203 VDD VSS sg13g2_decap_8
XFILLER_69_106 VDD VSS sg13g2_decap_8
XFILLER_3_861 VDD VSS sg13g2_decap_8
XFILLER_40_7 VDD VSS sg13g2_decap_8
XFILLER_97_459 VDD VSS sg13g2_decap_8
X_2250_ _2250_/RESET_B VSS VDD _2250_/D _2250_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_2_371 VDD VSS sg13g2_decap_8
XFILLER_78_640 VDD VSS sg13g2_fill_2
X_1201_ VDD _1201_/Y _1201_/A VSS sg13g2_inv_1
XIO_BOND_in_data_pads\[1\].in_data_pad in_data_PADs[1] bondpad_70x70
XFILLER_93_621 VDD VSS sg13g2_decap_8
X_2181_ _2181_/RESET_B VSS VDD _2181_/D _2181_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_77_161 VDD VSS sg13g2_decap_8
XFILLER_66_824 VDD VSS sg13g2_decap_8
XFILLER_93_665 VDD VSS sg13g2_decap_8
XFILLER_38_548 VDD VSS sg13g2_decap_8
XFILLER_81_849 VDD VSS sg13g2_decap_8
XFILLER_92_164 VDD VSS sg13g2_decap_8
XFILLER_65_378 VDD VSS sg13g2_decap_8
XFILLER_19_784 VDD VSS sg13g2_decap_8
XFILLER_80_348 VDD VSS sg13g2_decap_8
XFILLER_34_721 VDD VSS sg13g2_decap_8
XFILLER_18_294 VDD VSS sg13g2_decap_8
XFILLER_33_231 VDD VSS sg13g2_decap_8
XFILLER_22_938 VDD VSS sg13g2_decap_8
XFILLER_34_798 VDD VSS sg13g2_decap_8
X_1965_ _1961_/Y VDD _1966_/B VSS _1982_/A _1964_/D sg13g2_o21ai_1
XFILLER_21_448 VDD VSS sg13g2_decap_8
XFILLER_105_1043 VDD VSS sg13g2_decap_8
X_1896_ _1967_/A _1967_/B _1897_/A VDD VSS sg13g2_nor2b_1
X_2325__216 VDD VSS _2325_/RESET_B sg13g2_tiehi
XFILLER_108_49 VDD VSS sg13g2_decap_8
XFILLER_88_415 VDD VSS sg13g2_decap_8
XFILLER_0_308 VDD VSS sg13g2_decap_8
XFILLER_102_269 VDD VSS sg13g2_decap_8
XFILLER_64_1060 VDD VSS sg13g2_fill_1
XFILLER_25_1022 VDD VSS sg13g2_decap_8
XFILLER_29_504 VDD VSS sg13g2_decap_8
XFILLER_111_770 VDD VSS sg13g2_decap_8
XFILLER_56_312 VDD VSS sg13g2_decap_8
XFILLER_112_1036 VDD VSS sg13g2_decap_8
XFILLER_110_280 VDD VSS sg13g2_decap_8
XFILLER_68_183 VDD VSS sg13g2_decap_8
XFILLER_84_676 VDD VSS sg13g2_decap_8
XFILLER_71_315 VDD VSS sg13g2_decap_8
XFILLER_17_35 VDD VSS sg13g2_decap_8
XFILLER_44_529 VDD VSS sg13g2_decap_8
XFILLER_72_849 VDD VSS sg13g2_decap_4
XFILLER_37_581 VDD VSS sg13g2_decap_8
XFILLER_25_721 VDD VSS sg13g2_decap_8
XFILLER_80_860 VDD VSS sg13g2_fill_1
XFILLER_52_562 VDD VSS sg13g2_decap_8
XFILLER_52_540 VDD VSS sg13g2_decap_8
XFILLER_24_231 VDD VSS sg13g2_decap_8
XFILLER_40_746 VDD VSS sg13g2_decap_8
XFILLER_25_798 VDD VSS sg13g2_decap_8
XFILLER_13_938 VDD VSS sg13g2_decap_8
XFILLER_12_448 VDD VSS sg13g2_decap_8
XFILLER_33_56 VDD VSS sg13g2_decap_8
XFILLER_32_1015 VDD VSS sg13g2_decap_8
XFILLER_4_658 VDD VSS sg13g2_decap_8
XFILLER_3_168 VDD VSS sg13g2_decap_8
XFILLER_79_426 VDD VSS sg13g2_decap_8
XFILLER_0_875 VDD VSS sg13g2_decap_8
XFILLER_88_993 VDD VSS sg13g2_decap_8
XFILLER_48_835 VDD VSS sg13g2_decap_8
XFILLER_58_86 VDD VSS sg13g2_decap_8
XFILLER_75_665 VDD VSS sg13g2_decap_8
XFILLER_59_194 VDD VSS sg13g2_decap_8
XFILLER_47_345 VDD VSS sg13g2_decap_8
XFILLER_47_356 VDD VSS sg13g2_fill_2
XFILLER_35_518 VDD VSS sg13g2_decap_8
XFILLER_47_378 VDD VSS sg13g2_decap_8
XFILLER_74_63 VDD VSS sg13g2_decap_8
XFILLER_28_581 VDD VSS sg13g2_decap_8
XFILLER_62_337 VDD VSS sg13g2_decap_8
XFILLER_16_721 VDD VSS sg13g2_decap_8
XFILLER_90_668 VDD VSS sg13g2_decap_8
XFILLER_15_231 VDD VSS sg13g2_decap_8
XFILLER_71_893 VDD VSS sg13g2_decap_8
XFILLER_31_735 VDD VSS sg13g2_decap_8
XFILLER_16_798 VDD VSS sg13g2_decap_8
XFILLER_88_7 VDD VSS sg13g2_decap_8
XFILLER_30_245 VDD VSS sg13g2_decap_8
X_1750_ _1756_/B _1762_/A _1750_/A _1750_/Y VDD VSS sg13g2_nand3_1
XFILLER_90_84 VDD VSS sg13g2_decap_8
XFILLER_8_931 VDD VSS sg13g2_decap_8
XFILLER_7_441 VDD VSS sg13g2_decap_8
Xhold408 _2312_/Q VDD VSS _1680_/A sg13g2_dlygate4sd3_1
X_1681_ _1681_/A _1681_/B _2312_/D VDD VSS sg13g2_nor2_1
Xhold419 _2232_/Q VDD VSS _1422_/A sg13g2_dlygate4sd3_1
XFILLER_48_1044 VDD VSS sg13g2_decap_8
X_2302_ _2302_/RESET_B VSS VDD _2302_/D _2302_/Q _2369_/CLK sg13g2_dfrbpq_1
XFILLER_112_567 VDD VSS sg13g2_decap_8
XFILLER_97_256 VDD VSS sg13g2_decap_8
XFILLER_79_982 VDD VSS sg13g2_decap_8
X_2233_ _2233_/RESET_B VSS VDD _2233_/D _2233_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_66_610 VDD VSS sg13g2_fill_2
XFILLER_94_941 VDD VSS sg13g2_decap_8
X_2164_ _2164_/RESET_B VSS VDD _2164_/D _2164_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_39_857 VDD VSS sg13g2_decap_8
XFILLER_38_334 VDD VSS sg13g2_decap_8
XFILLER_26_518 VDD VSS sg13g2_decap_8
XFILLER_80_112 VDD VSS sg13g2_decap_4
XFILLER_19_581 VDD VSS sg13g2_decap_8
X_2095_ VDD _2095_/Y _2095_/A VSS sg13g2_inv_1
XFILLER_62_871 VDD VSS sg13g2_decap_8
XFILLER_0_1057 VDD VSS sg13g2_decap_4
XFILLER_80_178 VDD VSS sg13g2_decap_8
XFILLER_110_28 VDD VSS sg13g2_decap_8
XFILLER_34_595 VDD VSS sg13g2_decap_8
XFILLER_22_735 VDD VSS sg13g2_decap_8
XFILLER_55_1059 VDD VSS sg13g2_fill_2
XFILLER_21_245 VDD VSS sg13g2_decap_8
X_1948_ _1951_/A _1948_/A _1948_/B VDD VSS sg13g2_xnor2_1
XFILLER_9_91 VDD VSS sg13g2_decap_8
XFILLER_108_829 VDD VSS sg13g2_decap_8
X_1879_ _1887_/A _1879_/A _1879_/B VDD VSS sg13g2_xnor2_1
XFILLER_107_339 VDD VSS sg13g2_decap_8
XFILLER_89_713 VDD VSS sg13g2_decap_8
X_2329__193 VDD VSS _2329_/RESET_B sg13g2_tiehi
X_2184__172 VDD VSS _2184_/RESET_B sg13g2_tiehi
XFILLER_0_105 VDD VSS sg13g2_decap_8
XFILLER_77_919 VDD VSS sg13g2_decap_8
XFILLER_103_567 VDD VSS sg13g2_decap_8
XFILLER_76_429 VDD VSS sg13g2_decap_8
XFILLER_29_301 VDD VSS sg13g2_decap_8
XFILLER_57_632 VDD VSS sg13g2_decap_8
XFILLER_28_56 VDD VSS sg13g2_decap_8
XFILLER_56_131 VDD VSS sg13g2_decap_8
XFILLER_84_473 VDD VSS sg13g2_fill_2
XFILLER_17_518 VDD VSS sg13g2_decap_8
XFILLER_29_378 VDD VSS sg13g2_decap_8
XFILLER_44_315 VDD VSS sg13g2_decap_8
XFILLER_25_595 VDD VSS sg13g2_decap_8
XFILLER_13_735 VDD VSS sg13g2_decap_8
XFILLER_44_77 VDD VSS sg13g2_decap_8
XFILLER_40_543 VDD VSS sg13g2_decap_8
XFILLER_12_245 VDD VSS sg13g2_decap_8
XFILLER_9_728 VDD VSS sg13g2_decap_8
XFILLER_60_21 VDD VSS sg13g2_decap_4
XFILLER_8_238 VDD VSS sg13g2_decap_8
XFILLER_60_87 VDD VSS sg13g2_decap_8
XFILLER_5_945 VDD VSS sg13g2_decap_8
XFILLER_107_884 VDD VSS sg13g2_decap_8
XFILLER_109_70 VDD VSS sg13g2_decap_8
XFILLER_4_455 VDD VSS sg13g2_decap_8
XFILLER_5_49 VDD VSS sg13g2_decap_8
XFILLER_106_372 VDD VSS sg13g2_decap_8
XFILLER_48_610 VDD VSS sg13g2_decap_8
XFILLER_67_429 VDD VSS sg13g2_decap_8
XFILLER_0_672 VDD VSS sg13g2_decap_8
XFILLER_76_963 VDD VSS sg13g2_decap_8
XFILLER_75_440 VDD VSS sg13g2_decap_8
XFILLER_91_911 VDD VSS sg13g2_decap_4
Xclkbuf_2_3__f_clk clkbuf_leaf_9_clk/A clkbuf_0_clk/X VDD VSS sg13g2_buf_16
XFILLER_85_84 VDD VSS sg13g2_decap_8
XFILLER_48_687 VDD VSS sg13g2_decap_8
XFILLER_36_805 VDD VSS sg13g2_decap_8
XFILLER_91_933 VDD VSS sg13g2_decap_8
XFILLER_90_410 VDD VSS sg13g2_decap_8
XFILLER_63_635 VDD VSS sg13g2_decap_8
XFILLER_62_112 VDD VSS sg13g2_decap_8
XFILLER_35_315 VDD VSS sg13g2_decap_8
XFILLER_90_443 VDD VSS sg13g2_decap_8
XFILLER_62_134 VDD VSS sg13g2_decap_8
XFILLER_90_476 VDD VSS sg13g2_decap_8
XFILLER_44_893 VDD VSS sg13g2_decap_8
XFILLER_50_318 VDD VSS sg13g2_decap_8
X_2315__259 VDD VSS _2315_/RESET_B sg13g2_tiehi
XFILLER_71_690 VDD VSS sg13g2_decap_4
XFILLER_16_595 VDD VSS sg13g2_decap_8
XFILLER_31_532 VDD VSS sg13g2_decap_8
XFILLER_43_392 VDD VSS sg13g2_decap_8
X_1802_ VSS VDD _1801_/A _1801_/B _1802_/Y _1792_/Y sg13g2_a21oi_1
XFILLER_15_1043 VDD VSS sg13g2_decap_8
XFILLER_102_1013 VDD VSS sg13g2_decap_8
X_1733_ _1926_/B _2228_/Q _2236_/Q VDD VSS sg13g2_xnor2_1
X_1664_ _1670_/A _1664_/B _2304_/D VDD VSS sg13g2_nor2_1
XFILLER_98_532 VDD VSS sg13g2_decap_8
X_1595_ _1595_/A _1595_/B _1595_/Y VDD VSS sg13g2_nor2_1
XFILLER_59_908 VDD VSS sg13g2_decap_8
X_2361__279 VDD VSS _2361_/RESET_B sg13g2_tiehi
XFILLER_112_364 VDD VSS sg13g2_decap_8
XFILLER_105_28 VDD VSS sg13g2_decap_8
XFILLER_58_429 VDD VSS sg13g2_decap_8
X_2216_ _2216_/RESET_B VSS VDD _2216_/D _2216_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_85_259 VDD VSS sg13g2_decap_8
XFILLER_39_654 VDD VSS sg13g2_decap_8
XFILLER_82_900 VDD VSS sg13g2_decap_8
XFILLER_67_985 VDD VSS sg13g2_decap_8
XFILLER_22_1036 VDD VSS sg13g2_decap_8
XFILLER_27_805 VDD VSS sg13g2_decap_8
XFILLER_94_793 VDD VSS sg13g2_fill_2
XFILLER_93_270 VDD VSS sg13g2_decap_8
X_2147_ _2147_/A _2147_/B _2373_/D VDD VSS sg13g2_nor2_1
XFILLER_66_484 VDD VSS sg13g2_fill_2
XFILLER_26_315 VDD VSS sg13g2_decap_8
XFILLER_38_175 VDD VSS sg13g2_decap_8
XFILLER_82_977 VDD VSS sg13g2_decap_4
X_2078_ _2074_/Y VDD _2340_/D VSS _2076_/Y _2077_/Y sg13g2_o21ai_1
XFILLER_81_454 VDD VSS sg13g2_decap_8
XFILLER_54_668 VDD VSS sg13g2_fill_2
XFILLER_42_819 VDD VSS sg13g2_decap_8
XFILLER_35_882 VDD VSS sg13g2_decap_8
XFILLER_53_189 VDD VSS sg13g2_decap_8
XFILLER_41_329 VDD VSS sg13g2_decap_8
XFILLER_14_14 VDD VSS sg13g2_decap_8
XFILLER_22_532 VDD VSS sg13g2_decap_8
XFILLER_34_392 VDD VSS sg13g2_decap_8
XFILLER_10_749 VDD VSS sg13g2_decap_8
XFILLER_108_626 VDD VSS sg13g2_decap_8
XFILLER_30_35 VDD VSS sg13g2_decap_8
XFILLER_107_147 VDD VSS sg13g2_decap_8
XFILLER_104_865 VDD VSS sg13g2_decap_8
XFILLER_89_565 VDD VSS sg13g2_decap_8
XFILLER_103_320 VDD VSS sg13g2_decap_8
XFILLER_2_959 VDD VSS sg13g2_decap_8
XFILLER_7_1008 VDD VSS sg13g2_decap_8
XFILLER_77_716 VDD VSS sg13g2_decap_8
XFILLER_1_469 VDD VSS sg13g2_decap_8
XFILLER_103_397 VDD VSS sg13g2_decap_8
XFILLER_76_226 VDD VSS sg13g2_decap_8
XFILLER_39_77 VDD VSS sg13g2_decap_8
XFILLER_18_805 VDD VSS sg13g2_decap_8
XFILLER_72_421 VDD VSS sg13g2_decap_4
XFILLER_45_624 VDD VSS sg13g2_decap_8
XFILLER_17_315 VDD VSS sg13g2_decap_8
XFILLER_55_21 VDD VSS sg13g2_decap_8
XFILLER_29_175 VDD VSS sg13g2_decap_8
XFILLER_84_292 VDD VSS sg13g2_decap_8
XFILLER_60_605 VDD VSS sg13g2_decap_8
XFILLER_33_819 VDD VSS sg13g2_decap_8
XFILLER_44_134 VDD VSS sg13g2_decap_8
XFILLER_72_476 VDD VSS sg13g2_decap_8
XFILLER_38_1010 VDD VSS sg13g2_decap_8
XFILLER_26_882 VDD VSS sg13g2_decap_8
XFILLER_32_329 VDD VSS sg13g2_decap_8
XFILLER_53_690 VDD VSS sg13g2_decap_8
XFILLER_13_532 VDD VSS sg13g2_decap_8
XFILLER_25_392 VDD VSS sg13g2_decap_8
XFILLER_71_42 VDD VSS sg13g2_decap_8
XFILLER_41_874 VDD VSS sg13g2_decap_8
XFILLER_9_525 VDD VSS sg13g2_decap_8
XFILLER_40_384 VDD VSS sg13g2_decap_8
XFILLER_99_318 VDD VSS sg13g2_decap_8
XFILLER_5_742 VDD VSS sg13g2_decap_8
XFILLER_84_1030 VDD VSS sg13g2_decap_8
XFILLER_107_681 VDD VSS sg13g2_decap_8
XFILLER_4_252 VDD VSS sg13g2_decap_8
X_1380_ _1380_/Y _1380_/A _1389_/B VDD VSS sg13g2_nand2_1
XFILLER_45_1003 VDD VSS sg13g2_decap_8
XFILLER_110_802 VDD VSS sg13g2_decap_8
XFILLER_67_237 VDD VSS sg13g2_decap_8
XFILLER_110_879 VDD VSS sg13g2_decap_8
XFILLER_95_568 VDD VSS sg13g2_decap_8
XFILLER_83_719 VDD VSS sg13g2_decap_8
X_2001_ _2071_/B _2004_/B _2043_/S VDD VSS sg13g2_nor2b_1
XFILLER_49_974 VDD VSS sg13g2_decap_8
XFILLER_36_602 VDD VSS sg13g2_decap_8
XFILLER_48_451 VDD VSS sg13g2_decap_8
XFILLER_82_229 VDD VSS sg13g2_decap_8
XFILLER_64_944 VDD VSS sg13g2_decap_8
XFILLER_64_933 VDD VSS sg13g2_fill_2
XFILLER_64_922 VDD VSS sg13g2_decap_8
XFILLER_35_112 VDD VSS sg13g2_decap_8
XFILLER_91_752 VDD VSS sg13g2_decap_8
XFILLER_75_292 VDD VSS sg13g2_decap_8
XFILLER_51_605 VDD VSS sg13g2_decap_8
XFILLER_36_679 VDD VSS sg13g2_decap_8
XFILLER_24_819 VDD VSS sg13g2_decap_8
XFILLER_63_454 VDD VSS sg13g2_decap_8
XFILLER_17_882 VDD VSS sg13g2_decap_8
XFILLER_23_329 VDD VSS sg13g2_decap_8
XFILLER_35_189 VDD VSS sg13g2_decap_8
XFILLER_90_284 VDD VSS sg13g2_decap_4
XFILLER_44_690 VDD VSS sg13g2_decap_8
XFILLER_16_392 VDD VSS sg13g2_decap_8
XFILLER_91_1056 VDD VSS sg13g2_decap_4
XFILLER_52_1029 VDD VSS sg13g2_decap_8
XFILLER_52_1018 VDD VSS sg13g2_decap_4
XFILLER_32_896 VDD VSS sg13g2_decap_8
XFILLER_77_0 VDD VSS sg13g2_decap_8
X_1716_ _1716_/Y _1724_/S _1716_/B VDD VSS sg13g2_nand2_1
XFILLER_6_70 VDD VSS sg13g2_decap_8
X_1647_ _1674_/B _2328_/Q _2374_/Q _2343_/Q _2375_/Q _1677_/A _1647_/X VDD VSS sg13g2_mux4_1
XFILLER_86_524 VDD VSS sg13g2_decap_8
XFILLER_112_161 VDD VSS sg13g2_decap_8
X_1578_ VDD _1578_/Y _1578_/A VSS sg13g2_inv_1
XFILLER_58_215 VDD VSS sg13g2_decap_8
XFILLER_101_835 VDD VSS sg13g2_decap_8
XFILLER_86_535 VDD VSS sg13g2_fill_2
XFILLER_59_749 VDD VSS sg13g2_decap_8
XFILLER_58_248 VDD VSS sg13g2_decap_4
XFILLER_100_356 VDD VSS sg13g2_decap_8
XFILLER_27_602 VDD VSS sg13g2_decap_8
XFILLER_82_730 VDD VSS sg13g2_decap_8
XFILLER_73_229 VDD VSS sg13g2_decap_8
XFILLER_26_112 VDD VSS sg13g2_decap_8
XFILLER_55_966 VDD VSS sg13g2_decap_8
XFILLER_27_679 VDD VSS sg13g2_decap_8
XFILLER_54_432 VDD VSS sg13g2_decap_8
XFILLER_15_819 VDD VSS sg13g2_decap_8
XFILLER_109_1008 VDD VSS sg13g2_decap_8
XFILLER_82_785 VDD VSS sg13g2_decap_8
XFILLER_42_616 VDD VSS sg13g2_decap_8
XFILLER_14_329 VDD VSS sg13g2_decap_8
XFILLER_25_35 VDD VSS sg13g2_decap_8
XFILLER_26_189 VDD VSS sg13g2_decap_8
XFILLER_70_969 VDD VSS sg13g2_decap_8
XFILLER_81_284 VDD VSS sg13g2_decap_8
XFILLER_41_126 VDD VSS sg13g2_decap_8
XFILLER_50_671 VDD VSS sg13g2_decap_8
XFILLER_23_896 VDD VSS sg13g2_decap_8
XFILLER_109_924 VDD VSS sg13g2_decap_8
XFILLER_10_546 VDD VSS sg13g2_decap_8
XFILLER_41_56 VDD VSS sg13g2_decap_8
XFILLER_6_539 VDD VSS sg13g2_decap_8
XFILLER_108_478 VDD VSS sg13g2_decap_8
XFILLER_68_1047 VDD VSS sg13g2_decap_8
XFILLER_104_640 VDD VSS sg13g2_decap_8
XFILLER_2_756 VDD VSS sg13g2_decap_8
XFILLER_77_502 VDD VSS sg13g2_decap_8
XFILLER_1_266 VDD VSS sg13g2_decap_8
XFILLER_89_384 VDD VSS sg13g2_decap_8
XFILLER_103_161 VDD VSS sg13g2_decap_8
XFILLER_2_28 VDD VSS sg13g2_decap_8
XFILLER_77_579 VDD VSS sg13g2_decap_8
XFILLER_92_505 VDD VSS sg13g2_decap_8
XFILLER_46_911 VDD VSS sg13g2_decap_8
XFILLER_18_602 VDD VSS sg13g2_decap_8
XFILLER_66_42 VDD VSS sg13g2_decap_8
XFILLER_17_112 VDD VSS sg13g2_decap_8
XFILLER_45_421 VDD VSS sg13g2_decap_8
XFILLER_73_796 VDD VSS sg13g2_decap_8
XFILLER_33_616 VDD VSS sg13g2_decap_8
XFILLER_18_679 VDD VSS sg13g2_decap_8
XFILLER_45_476 VDD VSS sg13g2_decap_8
XFILLER_82_63 VDD VSS sg13g2_decap_8
XFILLER_61_969 VDD VSS sg13g2_fill_2
XFILLER_61_958 VDD VSS sg13g2_decap_8
XFILLER_60_424 VDD VSS sg13g2_fill_1
XFILLER_17_189 VDD VSS sg13g2_decap_8
XFILLER_32_126 VDD VSS sg13g2_decap_8
XFILLER_41_671 VDD VSS sg13g2_decap_8
XFILLER_9_322 VDD VSS sg13g2_decap_8
XFILLER_14_896 VDD VSS sg13g2_decap_8
XFILLER_70_7 VDD VSS sg13g2_decap_8
XFILLER_9_399 VDD VSS sg13g2_decap_8
XFILLER_12_1057 VDD VSS sg13g2_decap_4
XFILLER_108_990 VDD VSS sg13g2_decap_8
XFILLER_99_126 VDD VSS sg13g2_decap_8
X_1501_ _1501_/A _1501_/B _1518_/C VDD VSS sg13g2_nor2_1
X_1432_ _1433_/A _1429_/Y hold479/X _1429_/B _1370_/A VDD VSS sg13g2_a22oi_1
XFILLER_96_822 VDD VSS sg13g2_decap_8
XFILLER_95_321 VDD VSS sg13g2_decap_8
X_1363_ VDD _2210_/D _1363_/A VSS sg13g2_inv_1
XFILLER_110_676 VDD VSS sg13g2_decap_8
XFILLER_96_899 VDD VSS sg13g2_decap_8
X_1294_ _1294_/Y _1482_/B1 hold351/X _1482_/A2 _2341_/Q VDD VSS sg13g2_a22oi_1
XFILLER_68_579 VDD VSS sg13g2_decap_8
XFILLER_37_966 VDD VSS sg13g2_decap_8
XFILLER_48_281 VDD VSS sg13g2_decap_8
XFILLER_52_936 VDD VSS sg13g2_decap_8
XFILLER_64_774 VDD VSS sg13g2_decap_8
XFILLER_24_616 VDD VSS sg13g2_decap_8
XFILLER_63_262 VDD VSS sg13g2_decap_8
XFILLER_51_402 VDD VSS sg13g2_decap_4
XFILLER_36_476 VDD VSS sg13g2_decap_8
XFILLER_23_126 VDD VSS sg13g2_decap_8
XFILLER_32_693 VDD VSS sg13g2_decap_8
XFILLER_20_833 VDD VSS sg13g2_decap_8
XFILLER_106_916 VDD VSS sg13g2_decap_8
XFILLER_87_822 VDD VSS sg13g2_decap_8
XFILLER_86_321 VDD VSS sg13g2_decap_8
XFILLER_59_546 VDD VSS sg13g2_decap_8
XFILLER_101_643 VDD VSS sg13g2_fill_1
X_2300__111 VDD VSS _2300_/RESET_B sg13g2_tiehi
XFILLER_47_719 VDD VSS sg13g2_decap_8
XFILLER_98_1018 VDD VSS sg13g2_decap_8
XFILLER_86_398 VDD VSS sg13g2_decap_8
XFILLER_74_527 VDD VSS sg13g2_fill_1
XFILLER_100_164 VDD VSS sg13g2_fill_2
XFILLER_28_966 VDD VSS sg13g2_decap_8
XFILLER_55_741 VDD VSS sg13g2_decap_8
XFILLER_15_616 VDD VSS sg13g2_decap_8
XFILLER_36_56 VDD VSS sg13g2_decap_8
XFILLER_27_476 VDD VSS sg13g2_decap_8
XFILLER_43_947 VDD VSS sg13g2_decap_8
XFILLER_14_126 VDD VSS sg13g2_decap_8
XFILLER_70_766 VDD VSS sg13g2_decap_8
XFILLER_42_468 VDD VSS sg13g2_decap_8
XFILLER_23_693 VDD VSS sg13g2_decap_8
XFILLER_11_833 VDD VSS sg13g2_decap_8
XFILLER_35_1057 VDD VSS sg13g2_decap_4
XFILLER_10_343 VDD VSS sg13g2_decap_8
XFILLER_50_490 VDD VSS sg13g2_fill_2
XFILLER_109_721 VDD VSS sg13g2_decap_8
XFILLER_7_826 VDD VSS sg13g2_decap_8
XFILLER_6_336 VDD VSS sg13g2_decap_8
XFILLER_109_798 VDD VSS sg13g2_decap_8
XFILLER_108_264 VDD VSS sg13g2_fill_2
XFILLER_7_0 VDD VSS sg13g2_decap_8
XFILLER_81_1022 VDD VSS sg13g2_decap_8
XFILLER_2_553 VDD VSS sg13g2_decap_8
XFILLER_81_1055 VDD VSS sg13g2_decap_4
XFILLER_77_63 VDD VSS sg13g2_decap_8
XFILLER_78_888 VDD VSS sg13g2_decap_8
XFILLER_77_343 VDD VSS sg13g2_decap_8
XFILLER_93_825 VDD VSS sg13g2_decap_8
XFILLER_77_398 VDD VSS sg13g2_decap_8
XFILLER_19_966 VDD VSS sg13g2_decap_8
XFILLER_92_368 VDD VSS sg13g2_decap_8
XFILLER_93_84 VDD VSS sg13g2_decap_8
XFILLER_46_796 VDD VSS sg13g2_decap_8
XFILLER_34_903 VDD VSS sg13g2_decap_8
XFILLER_18_476 VDD VSS sg13g2_decap_8
XFILLER_45_262 VDD VSS sg13g2_decap_8
XFILLER_73_593 VDD VSS sg13g2_decap_8
XFILLER_60_221 VDD VSS sg13g2_decap_8
XFILLER_33_413 VDD VSS sg13g2_decap_8
X_1981_ VSS VDD _1982_/A _1982_/C _1995_/A _1982_/B sg13g2_a21oi_1
XFILLER_42_980 VDD VSS sg13g2_decap_8
XFILLER_14_693 VDD VSS sg13g2_decap_8
XFILLER_9_196 VDD VSS sg13g2_decap_8
XFILLER_96_630 VDD VSS sg13g2_decap_8
X_1415_ _1414_/Y VDD _2228_/D VSS _1370_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_111_952 VDD VSS sg13g2_decap_8
XFILLER_69_877 VDD VSS sg13g2_fill_1
XFILLER_95_140 VDD VSS sg13g2_decap_8
XFILLER_68_354 VDD VSS sg13g2_decap_8
X_1346_ _1366_/A _2266_/Q _2265_/Q _1409_/C _1346_/Y VDD VSS sg13g2_nor4_1
XFILLER_110_473 VDD VSS sg13g2_decap_8
Xout_data_pads\[5\].out_data_pad _2371_/Q IOVDD IOVSS out_data_PADs[5] VDD VSS sg13g2_IOPadOut30mA
X_1277_ VDD _2168_/D _1277_/A VSS sg13g2_inv_1
XFILLER_83_346 VDD VSS sg13g2_decap_8
XFILLER_3_1022 VDD VSS sg13g2_decap_8
XFILLER_64_571 VDD VSS sg13g2_decap_8
XFILLER_37_763 VDD VSS sg13g2_decap_8
XFILLER_25_903 VDD VSS sg13g2_decap_8
XFILLER_52_744 VDD VSS sg13g2_decap_8
XFILLER_19_1008 VDD VSS sg13g2_decap_8
XFILLER_24_413 VDD VSS sg13g2_decap_8
XFILLER_36_273 VDD VSS sg13g2_decap_8
XFILLER_40_928 VDD VSS sg13g2_decap_8
XFILLER_33_980 VDD VSS sg13g2_decap_8
XFILLER_51_298 VDD VSS sg13g2_decap_8
XFILLER_20_630 VDD VSS sg13g2_decap_8
XFILLER_22_14 VDD VSS sg13g2_decap_8
XFILLER_32_490 VDD VSS sg13g2_decap_8
XFILLER_106_713 VDD VSS sg13g2_decap_8
XFILLER_105_201 VDD VSS sg13g2_decap_8
XFILLER_105_256 VDD VSS sg13g2_decap_8
XFILLER_0_7 VDD VSS sg13g2_decap_8
XFILLER_87_630 VDD VSS sg13g2_decap_8
XFILLER_99_490 VDD VSS sg13g2_decap_8
XFILLER_102_963 VDD VSS sg13g2_decap_8
XFILLER_101_451 VDD VSS sg13g2_decap_8
XFILLER_87_696 VDD VSS sg13g2_decap_8
XFILLER_59_376 VDD VSS sg13g2_decap_8
XFILLER_47_516 VDD VSS sg13g2_decap_4
XFILLER_90_806 VDD VSS sg13g2_decap_8
XFILLER_75_869 VDD VSS sg13g2_decap_8
XFILLER_55_560 VDD VSS sg13g2_decap_8
XFILLER_28_763 VDD VSS sg13g2_decap_8
XFILLER_16_903 VDD VSS sg13g2_decap_8
X_2194__152 VDD VSS _2194_/RESET_B sg13g2_tiehi
XFILLER_43_744 VDD VSS sg13g2_decap_8
XFILLER_15_413 VDD VSS sg13g2_decap_8
XFILLER_63_21 VDD VSS sg13g2_decap_8
XFILLER_27_273 VDD VSS sg13g2_decap_8
XFILLER_70_563 VDD VSS sg13g2_decap_8
XFILLER_31_917 VDD VSS sg13g2_decap_8
XFILLER_24_980 VDD VSS sg13g2_decap_8
XFILLER_30_427 VDD VSS sg13g2_decap_8
XFILLER_42_287 VDD VSS sg13g2_decap_8
XFILLER_8_49 VDD VSS sg13g2_decap_8
XFILLER_11_630 VDD VSS sg13g2_decap_8
XFILLER_23_490 VDD VSS sg13g2_decap_8
XFILLER_10_140 VDD VSS sg13g2_decap_8
XFILLER_7_623 VDD VSS sg13g2_decap_8
XFILLER_6_133 VDD VSS sg13g2_decap_8
XFILLER_109_595 VDD VSS sg13g2_decap_8
XFILLER_12_91 VDD VSS sg13g2_decap_8
XFILLER_3_840 VDD VSS sg13g2_decap_8
XFILLER_98_917 VDD VSS sg13g2_decap_8
XFILLER_2_350 VDD VSS sg13g2_decap_8
XFILLER_112_749 VDD VSS sg13g2_decap_8
XFILLER_97_438 VDD VSS sg13g2_decap_8
XFILLER_88_84 VDD VSS sg13g2_decap_8
XFILLER_33_7 VDD VSS sg13g2_decap_8
XFILLER_78_652 VDD VSS sg13g2_decap_8
XFILLER_111_259 VDD VSS sg13g2_decap_8
XFILLER_77_140 VDD VSS sg13g2_decap_8
X_1200_ VDD _1200_/Y _1200_/A VSS sg13g2_inv_1
X_2180_ _2180_/RESET_B VSS VDD _2180_/D _2180_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_93_600 VDD VSS sg13g2_decap_8
XFILLER_65_313 VDD VSS sg13g2_decap_8
XFILLER_38_516 VDD VSS sg13g2_decap_4
XFILLER_65_335 VDD VSS sg13g2_fill_2
XFILLER_34_700 VDD VSS sg13g2_decap_8
XFILLER_19_763 VDD VSS sg13g2_decap_8
XFILLER_74_891 VDD VSS sg13g2_decap_8
XFILLER_80_327 VDD VSS sg13g2_decap_8
XFILLER_46_593 VDD VSS sg13g2_fill_1
XFILLER_18_273 VDD VSS sg13g2_decap_8
XFILLER_33_210 VDD VSS sg13g2_decap_8
XFILLER_22_917 VDD VSS sg13g2_decap_8
XFILLER_34_777 VDD VSS sg13g2_decap_8
XFILLER_15_980 VDD VSS sg13g2_decap_8
XFILLER_21_427 VDD VSS sg13g2_decap_8
XFILLER_33_287 VDD VSS sg13g2_decap_8
XFILLER_105_1022 VDD VSS sg13g2_decap_8
X_1964_ _1978_/A _1978_/B _1978_/C _1964_/D _1966_/A VDD VSS sg13g2_nor4_1
Xclkbuf_leaf_13_clk clkbuf_2_2__f_clk/X _2368_/CLK VDD VSS sg13g2_buf_8
XFILLER_14_490 VDD VSS sg13g2_decap_8
X_1895_ _1967_/B _1895_/A _1895_/B VDD VSS sg13g2_nand2_1
XFILLER_30_994 VDD VSS sg13g2_decap_8
XFILLER_108_28 VDD VSS sg13g2_decap_8
XFILLER_25_1001 VDD VSS sg13g2_decap_8
X_2260__231 VDD VSS _2260_/RESET_B sg13g2_tiehi
XFILLER_69_663 VDD VSS sg13g2_decap_8
XFILLER_112_1015 VDD VSS sg13g2_decap_8
XFILLER_69_685 VDD VSS sg13g2_decap_8
XFILLER_69_674 VDD VSS sg13g2_fill_1
XFILLER_57_814 VDD VSS sg13g2_fill_1
XFILLER_68_162 VDD VSS sg13g2_decap_8
XFILLER_84_655 VDD VSS sg13g2_decap_8
X_1329_ VDD _2194_/D _1329_/A VSS sg13g2_inv_1
XFILLER_96_493 VDD VSS sg13g2_decap_8
XFILLER_17_14 VDD VSS sg13g2_decap_8
XFILLER_72_828 VDD VSS sg13g2_decap_8
XFILLER_83_154 VDD VSS sg13g2_decap_8
XFILLER_37_560 VDD VSS sg13g2_decap_8
XFILLER_25_700 VDD VSS sg13g2_decap_8
XFILLER_44_508 VDD VSS sg13g2_decap_8
XFILLER_24_210 VDD VSS sg13g2_decap_8
XFILLER_80_850 VDD VSS sg13g2_fill_1
XFILLER_25_777 VDD VSS sg13g2_decap_8
XFILLER_13_917 VDD VSS sg13g2_decap_8
XFILLER_80_894 VDD VSS sg13g2_decap_8
XFILLER_40_725 VDD VSS sg13g2_decap_8
XFILLER_12_427 VDD VSS sg13g2_decap_8
XFILLER_24_287 VDD VSS sg13g2_decap_8
XFILLER_33_35 VDD VSS sg13g2_decap_8
XFILLER_71_1054 VDD VSS sg13g2_decap_8
XFILLER_21_994 VDD VSS sg13g2_decap_8
XFILLER_106_532 VDD VSS sg13g2_decap_8
XFILLER_4_637 VDD VSS sg13g2_decap_8
XFILLER_79_405 VDD VSS sg13g2_decap_8
XFILLER_3_147 VDD VSS sg13g2_decap_8
XFILLER_106_587 VDD VSS sg13g2_decap_8
XFILLER_58_21 VDD VSS sg13g2_fill_1
XFILLER_88_972 VDD VSS sg13g2_decap_8
XFILLER_0_854 VDD VSS sg13g2_decap_8
XFILLER_58_65 VDD VSS sg13g2_decap_8
XFILLER_94_419 VDD VSS sg13g2_decap_8
XFILLER_87_482 VDD VSS sg13g2_decap_8
XFILLER_48_814 VDD VSS sg13g2_decap_8
XFILLER_75_644 VDD VSS sg13g2_decap_8
XFILLER_87_493 VDD VSS sg13g2_fill_2
XFILLER_47_324 VDD VSS sg13g2_decap_8
XFILLER_74_154 VDD VSS sg13g2_decap_8
XFILLER_74_42 VDD VSS sg13g2_decap_8
XFILLER_63_839 VDD VSS sg13g2_decap_8
XFILLER_28_560 VDD VSS sg13g2_decap_8
XFILLER_16_700 VDD VSS sg13g2_decap_8
XFILLER_90_647 VDD VSS sg13g2_decap_8
XFILLER_62_316 VDD VSS sg13g2_decap_8
XFILLER_15_210 VDD VSS sg13g2_decap_8
XFILLER_71_861 VDD VSS sg13g2_fill_1
XFILLER_43_552 VDD VSS sg13g2_decap_8
XFILLER_16_777 VDD VSS sg13g2_decap_8
XFILLER_71_883 VDD VSS sg13g2_fill_1
XFILLER_43_563 VDD VSS sg13g2_fill_2
XFILLER_31_714 VDD VSS sg13g2_decap_8
XFILLER_15_287 VDD VSS sg13g2_decap_8
XFILLER_70_393 VDD VSS sg13g2_decap_8
XFILLER_90_63 VDD VSS sg13g2_decap_8
XFILLER_30_224 VDD VSS sg13g2_decap_8
XFILLER_8_910 VDD VSS sg13g2_decap_8
XFILLER_7_420 VDD VSS sg13g2_decap_8
XFILLER_12_994 VDD VSS sg13g2_decap_8
X_2224__92 VDD VSS _2224__92/L_HI sg13g2_tiehi
X_1680_ _1680_/B _1680_/A _1681_/B VDD VSS sg13g2_xor2_1
Xhold409 _2272_/Q VDD VSS _1260_/A sg13g2_dlygate4sd3_1
XFILLER_8_987 VDD VSS sg13g2_decap_8
XFILLER_109_392 VDD VSS sg13g2_decap_8
XFILLER_7_497 VDD VSS sg13g2_decap_8
XFILLER_48_1023 VDD VSS sg13g2_decap_8
X_2301_ _2301_/RESET_B VSS VDD _2301_/D _2301_/Q _2345_/CLK sg13g2_dfrbpq_1
XFILLER_98_725 VDD VSS sg13g2_decap_4
XFILLER_79_961 VDD VSS sg13g2_decap_8
XFILLER_112_546 VDD VSS sg13g2_decap_8
XFILLER_97_235 VDD VSS sg13g2_decap_8
XFILLER_94_920 VDD VSS sg13g2_decap_8
X_2232_ _2232_/RESET_B VSS VDD _2232_/D _2232_/Q clkload5/A sg13g2_dfrbpq_1
Xclkbuf_leaf_2_clk clkbuf_leaf_5_clk/A clkload5/A VDD VSS sg13g2_buf_8
XFILLER_39_836 VDD VSS sg13g2_decap_8
XFILLER_38_313 VDD VSS sg13g2_decap_8
X_2163_ _2163_/RESET_B VSS VDD _2163_/D _2163_/Q _2368_/CLK sg13g2_dfrbpq_1
XFILLER_94_997 VDD VSS sg13g2_decap_8
XFILLER_93_463 VDD VSS sg13g2_decap_8
XFILLER_19_560 VDD VSS sg13g2_decap_8
XFILLER_81_636 VDD VSS sg13g2_decap_8
XFILLER_47_880 VDD VSS sg13g2_decap_4
XFILLER_65_198 VDD VSS sg13g2_decap_8
XFILLER_53_338 VDD VSS sg13g2_decap_8
XFILLER_53_316 VDD VSS sg13g2_decap_8
XFILLER_53_327 VDD VSS sg13g2_fill_2
XFILLER_0_1036 VDD VSS sg13g2_decap_8
X_2094_ _2102_/B _2094_/B _2095_/A VDD VSS sg13g2_nor2_1
XFILLER_80_157 VDD VSS sg13g2_decap_8
XFILLER_62_850 VDD VSS sg13g2_decap_8
XFILLER_55_1038 VDD VSS sg13g2_decap_8
XFILLER_34_574 VDD VSS sg13g2_decap_8
XFILLER_22_714 VDD VSS sg13g2_decap_8
XFILLER_21_224 VDD VSS sg13g2_decap_8
XFILLER_9_70 VDD VSS sg13g2_decap_8
XFILLER_108_808 VDD VSS sg13g2_decap_8
X_1947_ VDD VSS _1984_/B _1945_/X _1984_/A _1985_/A _1978_/B _1985_/B sg13g2_a221oi_1
XFILLER_30_791 VDD VSS sg13g2_decap_8
X_1878_ _1879_/B _1878_/A _1878_/B VDD VSS sg13g2_xnor2_1
XFILLER_89_747 VDD VSS sg13g2_decap_8
XFILLER_88_213 VDD VSS sg13g2_decap_8
XFILLER_76_408 VDD VSS sg13g2_decap_8
XFILLER_57_611 VDD VSS sg13g2_decap_8
XFILLER_9_1050 VDD VSS sg13g2_decap_8
XFILLER_85_964 VDD VSS sg13g2_decap_8
XFILLER_28_35 VDD VSS sg13g2_decap_8
XFILLER_56_110 VDD VSS sg13g2_decap_8
XFILLER_84_452 VDD VSS sg13g2_decap_8
XFILLER_57_688 VDD VSS sg13g2_decap_8
XFILLER_45_828 VDD VSS sg13g2_decap_4
XFILLER_29_357 VDD VSS sg13g2_decap_8
XFILLER_84_496 VDD VSS sg13g2_decap_8
XFILLER_71_102 VDD VSS sg13g2_decap_4
XFILLER_38_891 VDD VSS sg13g2_decap_8
XFILLER_56_187 VDD VSS sg13g2_decap_8
XFILLER_53_894 VDD VSS sg13g2_decap_4
XFILLER_25_574 VDD VSS sg13g2_decap_8
XFILLER_13_714 VDD VSS sg13g2_decap_8
XFILLER_44_56 VDD VSS sg13g2_decap_8
XFILLER_52_382 VDD VSS sg13g2_decap_8
XFILLER_12_224 VDD VSS sg13g2_decap_8
XFILLER_9_707 VDD VSS sg13g2_decap_8
XFILLER_8_217 VDD VSS sg13g2_decap_8
XFILLER_100_84 VDD VSS sg13g2_decap_8
XFILLER_40_599 VDD VSS sg13g2_decap_8
XFILLER_21_791 VDD VSS sg13g2_decap_8
XFILLER_5_924 VDD VSS sg13g2_decap_8
XFILLER_60_66 VDD VSS sg13g2_decap_8
XFILLER_4_434 VDD VSS sg13g2_decap_8
XFILLER_5_28 VDD VSS sg13g2_decap_8
XFILLER_107_863 VDD VSS sg13g2_decap_8
XFILLER_106_340 VDD VSS sg13g2_decap_4
XFILLER_107_0 VDD VSS sg13g2_decap_8
XFILLER_79_224 VDD VSS sg13g2_decap_4
XFILLER_69_42 VDD VSS sg13g2_decap_8
XFILLER_79_257 VDD VSS sg13g2_fill_1
XFILLER_67_408 VDD VSS sg13g2_decap_8
XFILLER_0_651 VDD VSS sg13g2_decap_8
XFILLER_87_290 VDD VSS sg13g2_decap_8
XFILLER_85_63 VDD VSS sg13g2_decap_8
XFILLER_63_614 VDD VSS sg13g2_decap_8
XFILLER_48_666 VDD VSS sg13g2_decap_8
XFILLER_47_132 VDD VSS sg13g2_decap_8
XFILLER_78_1049 VDD VSS sg13g2_decap_8
XFILLER_47_198 VDD VSS sg13g2_decap_8
XFILLER_44_872 VDD VSS sg13g2_decap_8
XFILLER_16_574 VDD VSS sg13g2_decap_8
XFILLER_31_511 VDD VSS sg13g2_decap_8
XFILLER_43_371 VDD VSS sg13g2_decap_8
X_1801_ _1801_/Y _1801_/A _1801_/B VDD VSS sg13g2_nand2_1
XFILLER_15_1022 VDD VSS sg13g2_decap_8
XFILLER_31_588 VDD VSS sg13g2_decap_8
XFILLER_12_791 VDD VSS sg13g2_decap_8
X_1732_ _2236_/Q _2228_/Q _1732_/Y VDD VSS sg13g2_nor2b_1
X_1663_ _1663_/Y _1646_/Y _1662_/X hold427/X _1189_/Y VDD VSS sg13g2_a22oi_1
XFILLER_8_784 VDD VSS sg13g2_decap_8
XFILLER_7_294 VDD VSS sg13g2_decap_8
XFILLER_98_511 VDD VSS sg13g2_decap_8
X_1594_ _1595_/B _1594_/A _1594_/B VDD VSS sg13g2_xnor2_1
XIO_FILL_IO_EAST_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_112_343 VDD VSS sg13g2_decap_8
XFILLER_98_588 VDD VSS sg13g2_decap_8
XFILLER_86_739 VDD VSS sg13g2_decap_8
XFILLER_22_0 VDD VSS sg13g2_decap_8
XFILLER_100_538 VDD VSS sg13g2_decap_8
X_2215_ _2215_/RESET_B VSS VDD _2215_/D _2215_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_85_238 VDD VSS sg13g2_decap_8
XFILLER_22_1015 VDD VSS sg13g2_decap_8
XFILLER_39_633 VDD VSS sg13g2_decap_8
XFILLER_94_772 VDD VSS sg13g2_decap_8
XFILLER_67_964 VDD VSS sg13g2_decap_8
XFILLER_66_463 VDD VSS sg13g2_decap_8
XFILLER_38_154 VDD VSS sg13g2_decap_8
XFILLER_82_956 VDD VSS sg13g2_decap_8
X_2146_ _1688_/B VDD _2147_/B VSS hold564/X _1259_/A sg13g2_o21ai_1
XFILLER_54_647 VDD VSS sg13g2_decap_8
X_2077_ _2077_/A _2089_/S _2077_/Y VDD VSS sg13g2_nor2b_1
XFILLER_81_433 VDD VSS sg13g2_decap_8
XFILLER_53_146 VDD VSS sg13g2_decap_4
XFILLER_35_861 VDD VSS sg13g2_decap_8
XFILLER_41_308 VDD VSS sg13g2_decap_8
XFILLER_22_511 VDD VSS sg13g2_decap_8
XFILLER_34_371 VDD VSS sg13g2_decap_8
XFILLER_22_588 VDD VSS sg13g2_decap_8
XFILLER_10_728 VDD VSS sg13g2_decap_8
XFILLER_108_605 VDD VSS sg13g2_decap_8
XFILLER_30_14 VDD VSS sg13g2_decap_8
XFILLER_107_126 VDD VSS sg13g2_decap_8
XFILLER_100_7 VDD VSS sg13g2_decap_8
XFILLER_2_938 VDD VSS sg13g2_decap_8
XFILLER_89_544 VDD VSS sg13g2_decap_8
XFILLER_1_448 VDD VSS sg13g2_decap_8
XFILLER_103_376 VDD VSS sg13g2_decap_8
XFILLER_39_56 VDD VSS sg13g2_decap_8
XFILLER_49_419 VDD VSS sg13g2_decap_8
XFILLER_73_901 VDD VSS sg13g2_decap_8
XFILLER_29_154 VDD VSS sg13g2_decap_8
XFILLER_84_271 VDD VSS sg13g2_decap_8
XFILLER_72_400 VDD VSS sg13g2_decap_8
XFILLER_73_967 VDD VSS sg13g2_decap_8
XFILLER_72_455 VDD VSS sg13g2_decap_8
XFILLER_45_647 VDD VSS sg13g2_decap_4
XFILLER_77_1060 VDD VSS sg13g2_fill_1
XFILLER_26_861 VDD VSS sg13g2_decap_8
XFILLER_55_88 VDD VSS sg13g2_decap_8
XFILLER_32_308 VDD VSS sg13g2_decap_8
XFILLER_71_21 VDD VSS sg13g2_decap_8
XFILLER_41_853 VDD VSS sg13g2_decap_8
XFILLER_13_511 VDD VSS sg13g2_decap_8
XFILLER_25_371 VDD VSS sg13g2_decap_8
XFILLER_9_504 VDD VSS sg13g2_decap_8
XFILLER_40_363 VDD VSS sg13g2_decap_8
XFILLER_13_588 VDD VSS sg13g2_decap_8
XFILLER_5_721 VDD VSS sg13g2_decap_8
XFILLER_4_231 VDD VSS sg13g2_decap_8
XFILLER_107_660 VDD VSS sg13g2_decap_8
XFILLER_5_798 VDD VSS sg13g2_decap_8
XFILLER_20_91 VDD VSS sg13g2_decap_8
XFILLER_95_503 VDD VSS sg13g2_decap_8
XFILLER_45_1059 VDD VSS sg13g2_fill_2
XFILLER_110_858 VDD VSS sg13g2_decap_8
XFILLER_95_536 VDD VSS sg13g2_decap_8
XFILLER_96_84 VDD VSS sg13g2_decap_8
XFILLER_49_931 VDD VSS sg13g2_decap_8
XFILLER_67_216 VDD VSS sg13g2_decap_8
X_2000_ _2000_/B _2000_/C _2000_/A _2004_/B VDD VSS sg13g2_nand3_1
XFILLER_82_208 VDD VSS sg13g2_decap_8
XFILLER_64_901 VDD VSS sg13g2_decap_8
XFILLER_48_430 VDD VSS sg13g2_decap_8
XFILLER_91_731 VDD VSS sg13g2_decap_8
XFILLER_76_783 VDD VSS sg13g2_decap_8
XFILLER_75_271 VDD VSS sg13g2_decap_8
XFILLER_48_496 VDD VSS sg13g2_decap_8
XFILLER_36_658 VDD VSS sg13g2_decap_8
XFILLER_63_433 VDD VSS sg13g2_decap_8
XFILLER_90_263 VDD VSS sg13g2_decap_8
XFILLER_17_861 VDD VSS sg13g2_decap_8
XFILLER_23_308 VDD VSS sg13g2_decap_8
XFILLER_35_168 VDD VSS sg13g2_decap_8
XFILLER_91_1035 VDD VSS sg13g2_decap_8
XFILLER_16_371 VDD VSS sg13g2_decap_8
XFILLER_50_127 VDD VSS sg13g2_decap_8
XFILLER_32_875 VDD VSS sg13g2_decap_8
XFILLER_31_385 VDD VSS sg13g2_decap_8
X_1715_ _1716_/B _1715_/A _1719_/B VDD VSS sg13g2_xnor2_1
XFILLER_8_581 VDD VSS sg13g2_decap_8
X_2285__167 VDD VSS _2285_/RESET_B sg13g2_tiehi
X_1646_ _2312_/Q _1671_/B _1646_/Y VDD VSS sg13g2_nor2_1
XFILLER_99_864 VDD VSS sg13g2_fill_2
X_1577_ _1577_/S0 _2242_/Q _2234_/Q _2226_/Q _2218_/Q _2287_/Q _1578_/A VDD VSS sg13g2_mux4_1
XFILLER_101_814 VDD VSS sg13g2_decap_8
XFILLER_112_140 VDD VSS sg13g2_decap_8
XFILLER_59_728 VDD VSS sg13g2_decap_8
XFILLER_101_858 VDD VSS sg13g2_decap_8
XFILLER_101_869 VDD VSS sg13g2_fill_1
XFILLER_74_709 VDD VSS sg13g2_decap_8
XFILLER_73_208 VDD VSS sg13g2_decap_8
XFILLER_94_580 VDD VSS sg13g2_decap_8
XFILLER_66_260 VDD VSS sg13g2_fill_1
XFILLER_66_271 VDD VSS sg13g2_decap_8
XFILLER_54_411 VDD VSS sg13g2_decap_8
XFILLER_39_485 VDD VSS sg13g2_decap_8
X_2129_ VDD VSS _2124_/B _2120_/A _2128_/X hold345/X _2131_/A _2124_/Y sg13g2_a221oi_1
XFILLER_27_658 VDD VSS sg13g2_decap_8
XFILLER_81_263 VDD VSS sg13g2_decap_8
XFILLER_54_488 VDD VSS sg13g2_decap_8
XFILLER_14_308 VDD VSS sg13g2_decap_8
XFILLER_25_14 VDD VSS sg13g2_decap_8
XFILLER_41_105 VDD VSS sg13g2_decap_8
XFILLER_26_168 VDD VSS sg13g2_decap_8
XFILLER_70_948 VDD VSS sg13g2_decap_8
XFILLER_50_650 VDD VSS sg13g2_decap_8
XFILLER_23_875 VDD VSS sg13g2_decap_8
XFILLER_10_525 VDD VSS sg13g2_decap_8
XFILLER_22_385 VDD VSS sg13g2_decap_8
XFILLER_109_903 VDD VSS sg13g2_decap_8
XFILLER_6_518 VDD VSS sg13g2_decap_8
XFILLER_41_35 VDD VSS sg13g2_decap_8
XFILLER_108_457 VDD VSS sg13g2_decap_8
Xhold570 _2266_/Q VDD VSS _1192_/A sg13g2_dlygate4sd3_1
XFILLER_2_735 VDD VSS sg13g2_decap_8
XFILLER_89_363 VDD VSS sg13g2_decap_4
XFILLER_103_140 VDD VSS sg13g2_decap_8
XFILLER_1_245 VDD VSS sg13g2_decap_8
XFILLER_104_696 VDD VSS sg13g2_decap_8
XFILLER_77_558 VDD VSS sg13g2_decap_8
X_2240__262 VDD VSS _2240_/RESET_B sg13g2_tiehi
XFILLER_66_21 VDD VSS sg13g2_decap_8
XFILLER_64_219 VDD VSS sg13g2_decap_8
XFILLER_18_658 VDD VSS sg13g2_decap_8
XFILLER_66_98 VDD VSS sg13g2_decap_8
XFILLER_45_455 VDD VSS sg13g2_decap_8
XFILLER_75_1019 VDD VSS sg13g2_fill_1
XFILLER_46_989 VDD VSS sg13g2_decap_8
XFILLER_17_168 VDD VSS sg13g2_decap_8
XFILLER_32_105 VDD VSS sg13g2_decap_8
XFILLER_82_42 VDD VSS sg13g2_decap_8
XFILLER_41_650 VDD VSS sg13g2_decap_8
XFILLER_9_301 VDD VSS sg13g2_decap_8
XFILLER_14_875 VDD VSS sg13g2_decap_8
XFILLER_13_385 VDD VSS sg13g2_decap_8
XFILLER_15_91 VDD VSS sg13g2_decap_8
XFILLER_51_1052 VDD VSS sg13g2_decap_8
XFILLER_40_182 VDD VSS sg13g2_decap_8
XFILLER_9_378 VDD VSS sg13g2_decap_8
XFILLER_12_1036 VDD VSS sg13g2_decap_8
XFILLER_63_7 VDD VSS sg13g2_decap_8
XFILLER_99_105 VDD VSS sg13g2_decap_8
X_1500_ _1500_/A _1500_/B _2355_/Q _1500_/D _1518_/B VDD VSS sg13g2_nor4_1
X_1431_ VDD _2235_/D _1431_/A VSS sg13g2_inv_1
XFILLER_5_595 VDD VSS sg13g2_decap_8
XFILLER_95_300 VDD VSS sg13g2_decap_8
X_1362_ _1363_/A _1347_/Y hold449/X _1347_/B _1388_/A VDD VSS sg13g2_a22oi_1
XFILLER_110_655 VDD VSS sg13g2_decap_8
XFILLER_96_878 VDD VSS sg13g2_decap_8
X_1293_ VDD _2176_/D _1293_/A VSS sg13g2_inv_1
XFILLER_68_558 VDD VSS sg13g2_decap_8
XFILLER_95_399 VDD VSS sg13g2_decap_8
XFILLER_49_783 VDD VSS sg13g2_decap_8
XFILLER_48_260 VDD VSS sg13g2_decap_8
XFILLER_37_945 VDD VSS sg13g2_decap_8
XFILLER_64_753 VDD VSS sg13g2_decap_8
XFILLER_52_915 VDD VSS sg13g2_decap_8
XFILLER_36_455 VDD VSS sg13g2_decap_8
XFILLER_51_436 VDD VSS sg13g2_decap_8
XFILLER_23_105 VDD VSS sg13g2_decap_8
XFILLER_51_458 VDD VSS sg13g2_fill_1
XFILLER_108_1053 VDD VSS sg13g2_decap_8
XFILLER_60_970 VDD VSS sg13g2_decap_8
XFILLER_32_672 VDD VSS sg13g2_decap_8
XFILLER_20_812 VDD VSS sg13g2_decap_8
XFILLER_31_182 VDD VSS sg13g2_decap_8
XFILLER_20_889 VDD VSS sg13g2_decap_8
XFILLER_11_49 VDD VSS sg13g2_decap_8
XFILLER_105_449 VDD VSS sg13g2_decap_8
X_1629_ _1630_/B _1629_/A _1633_/B VDD VSS sg13g2_xnor2_1
XFILLER_87_801 VDD VSS sg13g2_decap_8
XFILLER_28_1043 VDD VSS sg13g2_decap_8
XFILLER_101_622 VDD VSS sg13g2_decap_8
XFILLER_99_694 VDD VSS sg13g2_decap_8
XFILLER_59_525 VDD VSS sg13g2_decap_8
XFILLER_98_1008 VDD VSS sg13g2_decap_4
XFILLER_101_655 VDD VSS sg13g2_fill_2
XFILLER_87_878 VDD VSS sg13g2_decap_8
XFILLER_101_699 VDD VSS sg13g2_decap_8
XFILLER_86_377 VDD VSS sg13g2_decap_8
XFILLER_100_154 VDD VSS sg13g2_fill_2
XFILLER_55_720 VDD VSS sg13g2_decap_8
XFILLER_100_198 VDD VSS sg13g2_decap_4
XFILLER_28_945 VDD VSS sg13g2_decap_8
XFILLER_36_35 VDD VSS sg13g2_decap_8
XFILLER_43_926 VDD VSS sg13g2_decap_8
X_2374__257 VDD VSS _2374_/RESET_B sg13g2_tiehi
XFILLER_54_252 VDD VSS sg13g2_decap_4
XFILLER_27_455 VDD VSS sg13g2_decap_8
XFILLER_82_583 VDD VSS sg13g2_decap_8
XFILLER_70_745 VDD VSS sg13g2_decap_8
XFILLER_55_797 VDD VSS sg13g2_decap_8
XFILLER_54_285 VDD VSS sg13g2_decap_8
XFILLER_14_105 VDD VSS sg13g2_decap_8
XFILLER_74_1052 VDD VSS sg13g2_decap_8
XFILLER_30_609 VDD VSS sg13g2_decap_8
XFILLER_42_447 VDD VSS sg13g2_decap_8
XFILLER_35_1036 VDD VSS sg13g2_decap_8
XFILLER_23_672 VDD VSS sg13g2_decap_8
XFILLER_11_812 VDD VSS sg13g2_decap_8
XFILLER_109_700 VDD VSS sg13g2_decap_8
XFILLER_10_322 VDD VSS sg13g2_decap_8
XFILLER_7_805 VDD VSS sg13g2_decap_8
XFILLER_52_89 VDD VSS sg13g2_decap_8
XFILLER_22_182 VDD VSS sg13g2_decap_8
XFILLER_6_315 VDD VSS sg13g2_decap_8
XFILLER_11_889 VDD VSS sg13g2_decap_8
XFILLER_108_243 VDD VSS sg13g2_decap_8
XFILLER_10_399 VDD VSS sg13g2_decap_8
XFILLER_109_777 VDD VSS sg13g2_decap_8
XFILLER_108_298 VDD VSS sg13g2_decap_4
XFILLER_2_532 VDD VSS sg13g2_decap_8
XFILLER_105_994 VDD VSS sg13g2_decap_8
XFILLER_81_1034 VDD VSS sg13g2_decap_8
XFILLER_78_845 VDD VSS sg13g2_fill_2
XFILLER_78_834 VDD VSS sg13g2_decap_8
XFILLER_77_322 VDD VSS sg13g2_decap_8
XFILLER_96_119 VDD VSS sg13g2_decap_8
XFILLER_77_42 VDD VSS sg13g2_decap_8
XFILLER_93_804 VDD VSS sg13g2_decap_8
XFILLER_89_193 VDD VSS sg13g2_decap_8
XFILLER_42_1029 VDD VSS sg13g2_decap_8
XFILLER_38_709 VDD VSS sg13g2_decap_8
XFILLER_77_377 VDD VSS sg13g2_decap_8
XFILLER_93_859 VDD VSS sg13g2_decap_8
XFILLER_92_347 VDD VSS sg13g2_decap_8
XFILLER_19_945 VDD VSS sg13g2_decap_8
XFILLER_80_509 VDD VSS sg13g2_decap_8
XFILLER_93_63 VDD VSS sg13g2_decap_8
XFILLER_46_775 VDD VSS sg13g2_decap_8
XFILLER_18_455 VDD VSS sg13g2_decap_8
XFILLER_34_959 VDD VSS sg13g2_decap_8
XFILLER_60_200 VDD VSS sg13g2_decap_8
X_1980_ _2000_/B _1982_/C _1980_/B VDD VSS sg13g2_nand2_1
XFILLER_21_609 VDD VSS sg13g2_decap_8
XFILLER_33_469 VDD VSS sg13g2_decap_8
XFILLER_60_277 VDD VSS sg13g2_decap_8
XFILLER_20_119 VDD VSS sg13g2_decap_8
XFILLER_14_672 VDD VSS sg13g2_decap_8
XFILLER_13_182 VDD VSS sg13g2_decap_8
XFILLER_9_175 VDD VSS sg13g2_decap_8
XFILLER_6_882 VDD VSS sg13g2_decap_8
XFILLER_5_392 VDD VSS sg13g2_decap_8
XFILLER_111_931 VDD VSS sg13g2_decap_8
XFILLER_69_823 VDD VSS sg13g2_decap_8
X_1414_ _1414_/Y _1414_/A _1426_/B VDD VSS sg13g2_nand2_1
X_1345_ VDD _2202_/D _1345_/A VSS sg13g2_inv_1
XFILLER_68_333 VDD VSS sg13g2_decap_8
XFILLER_96_686 VDD VSS sg13g2_decap_8
XFILLER_110_452 VDD VSS sg13g2_decap_8
XFILLER_68_399 VDD VSS sg13g2_decap_8
XFILLER_3_1001 VDD VSS sg13g2_decap_8
X_1276_ _1276_/Y _1338_/B1 hold302/X _1338_/A2 _2318_/Q VDD VSS sg13g2_a22oi_1
XFILLER_95_196 VDD VSS sg13g2_decap_8
XFILLER_83_358 VDD VSS sg13g2_fill_2
XFILLER_37_742 VDD VSS sg13g2_decap_8
XFILLER_71_509 VDD VSS sg13g2_decap_8
XFILLER_64_550 VDD VSS sg13g2_decap_8
XFILLER_52_712 VDD VSS sg13g2_decap_8
XFILLER_36_252 VDD VSS sg13g2_decap_8
XFILLER_25_959 VDD VSS sg13g2_decap_8
XFILLER_52_734 VDD VSS sg13g2_decap_4
XFILLER_40_907 VDD VSS sg13g2_decap_8
XFILLER_12_609 VDD VSS sg13g2_decap_8
XFILLER_24_469 VDD VSS sg13g2_decap_8
XFILLER_51_244 VDD VSS sg13g2_decap_8
XFILLER_11_119 VDD VSS sg13g2_decap_8
XFILLER_20_686 VDD VSS sg13g2_decap_8
XFILLER_4_819 VDD VSS sg13g2_decap_8
XFILLER_105_235 VDD VSS sg13g2_decap_8
XFILLER_3_329 VDD VSS sg13g2_decap_8
XFILLER_106_769 VDD VSS sg13g2_decap_8
XFILLER_65_1029 VDD VSS sg13g2_decap_8
XFILLER_102_920 VDD VSS sg13g2_fill_2
XFILLER_78_119 VDD VSS sg13g2_decap_8
XFILLER_102_942 VDD VSS sg13g2_decap_8
XFILLER_101_430 VDD VSS sg13g2_decap_8
XFILLER_59_355 VDD VSS sg13g2_decap_8
XFILLER_87_675 VDD VSS sg13g2_decap_8
XFILLER_74_314 VDD VSS sg13g2_decap_8
XFILLER_75_848 VDD VSS sg13g2_decap_8
XFILLER_86_185 VDD VSS sg13g2_decap_8
XFILLER_28_742 VDD VSS sg13g2_decap_8
XFILLER_47_56 VDD VSS sg13g2_decap_8
XFILLER_47_539 VDD VSS sg13g2_fill_2
XFILLER_27_252 VDD VSS sg13g2_decap_8
XFILLER_83_892 VDD VSS sg13g2_decap_8
XFILLER_103_84 VDD VSS sg13g2_decap_8
XFILLER_43_723 VDD VSS sg13g2_decap_8
XFILLER_16_959 VDD VSS sg13g2_decap_8
XFILLER_70_542 VDD VSS sg13g2_decap_8
XFILLER_15_469 VDD VSS sg13g2_decap_8
Xout_valid_pad _2273_/Q IOVDD IOVSS out_valid_PAD VDD VSS sg13g2_IOPadOut30mA
XFILLER_30_406 VDD VSS sg13g2_decap_8
XFILLER_42_266 VDD VSS sg13g2_decap_8
XFILLER_8_28 VDD VSS sg13g2_decap_8
XFILLER_7_602 VDD VSS sg13g2_decap_8
XFILLER_6_112 VDD VSS sg13g2_decap_8
XFILLER_11_686 VDD VSS sg13g2_decap_8
XFILLER_109_574 VDD VSS sg13g2_decap_8
XFILLER_10_196 VDD VSS sg13g2_decap_8
XFILLER_12_70 VDD VSS sg13g2_decap_8
XFILLER_7_679 VDD VSS sg13g2_decap_8
XFILLER_98_907 VDD VSS sg13g2_fill_1
XFILLER_6_189 VDD VSS sg13g2_decap_8
XFILLER_88_63 VDD VSS sg13g2_decap_8
XFILLER_112_728 VDD VSS sg13g2_decap_8
XFILLER_105_791 VDD VSS sg13g2_decap_8
XFILLER_3_896 VDD VSS sg13g2_decap_8
XFILLER_111_238 VDD VSS sg13g2_decap_8
XFILLER_26_7 VDD VSS sg13g2_decap_8
XFILLER_78_697 VDD VSS sg13g2_decap_8
XFILLER_93_656 VDD VSS sg13g2_fill_1
XFILLER_77_196 VDD VSS sg13g2_decap_8
XFILLER_19_742 VDD VSS sg13g2_decap_8
XFILLER_80_306 VDD VSS sg13g2_decap_8
XFILLER_18_252 VDD VSS sg13g2_decap_8
XFILLER_92_199 VDD VSS sg13g2_decap_8
XFILLER_34_756 VDD VSS sg13g2_decap_8
XFILLER_61_597 VDD VSS sg13g2_decap_8
XFILLER_21_406 VDD VSS sg13g2_decap_8
XFILLER_33_266 VDD VSS sg13g2_decap_8
XFILLER_105_1001 VDD VSS sg13g2_decap_8
X_1963_ VDD _1964_/D _1982_/B VSS sg13g2_inv_1
X_1894_ _1895_/B _1960_/A _1960_/B VDD VSS sg13g2_nand2_1
XFILLER_30_973 VDD VSS sg13g2_decap_8
XFILLER_88_1007 VDD VSS sg13g2_decap_8
XFILLER_88_1018 VDD VSS sg13g2_fill_2
XIO_FILL_IO_SOUTH_7_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_52_0 VDD VSS sg13g2_decap_8
XFILLER_89_929 VDD VSS sg13g2_decap_8
XFILLER_102_205 VDD VSS sg13g2_decap_4
XFILLER_69_642 VDD VSS sg13g2_decap_8
XFILLER_97_984 VDD VSS sg13g2_decap_8
XFILLER_84_601 VDD VSS sg13g2_fill_1
XFILLER_25_1057 VDD VSS sg13g2_decap_4
XFILLER_84_634 VDD VSS sg13g2_decap_8
X_1328_ _1328_/Y _1344_/B1 hold381/X _1344_/A2 _2327_/Q VDD VSS sg13g2_a22oi_1
XFILLER_83_133 VDD VSS sg13g2_decap_4
XFILLER_56_347 VDD VSS sg13g2_decap_8
XFILLER_29_539 VDD VSS sg13g2_decap_8
X_1259_ _2273_/Q _1259_/C _1259_/A _1514_/A VDD VSS sg13g2_nand3_1
XFILLER_83_199 VDD VSS sg13g2_decap_8
XFILLER_65_881 VDD VSS sg13g2_decap_8
XFILLER_25_756 VDD VSS sg13g2_decap_8
XFILLER_40_704 VDD VSS sg13g2_decap_8
XFILLER_12_406 VDD VSS sg13g2_decap_8
XFILLER_33_14 VDD VSS sg13g2_decap_8
XFILLER_24_266 VDD VSS sg13g2_decap_8
XFILLER_71_1033 VDD VSS sg13g2_decap_8
XFILLER_21_973 VDD VSS sg13g2_decap_8
XFILLER_20_483 VDD VSS sg13g2_decap_8
XFILLER_4_616 VDD VSS sg13g2_decap_8
XFILLER_106_511 VDD VSS sg13g2_decap_8
XFILLER_3_126 VDD VSS sg13g2_decap_8
XFILLER_106_566 VDD VSS sg13g2_decap_8
XFILLER_0_833 VDD VSS sg13g2_decap_8
XFILLER_59_141 VDD VSS sg13g2_decap_4
XFILLER_59_152 VDD VSS sg13g2_fill_2
XFILLER_75_623 VDD VSS sg13g2_decap_8
XFILLER_47_314 VDD VSS sg13g2_fill_1
XFILLER_90_615 VDD VSS sg13g2_decap_8
XFILLER_74_133 VDD VSS sg13g2_decap_8
XFILLER_74_21 VDD VSS sg13g2_decap_8
XFILLER_63_818 VDD VSS sg13g2_decap_8
XFILLER_56_892 VDD VSS sg13g2_decap_8
XFILLER_71_840 VDD VSS sg13g2_decap_8
XFILLER_74_98 VDD VSS sg13g2_decap_8
XFILLER_16_756 VDD VSS sg13g2_decap_8
XFILLER_70_372 VDD VSS sg13g2_decap_8
XFILLER_15_266 VDD VSS sg13g2_decap_8
XFILLER_30_203 VDD VSS sg13g2_decap_8
XFILLER_90_42 VDD VSS sg13g2_decap_8
XFILLER_43_597 VDD VSS sg13g2_decap_8
XFILLER_12_973 VDD VSS sg13g2_decap_8
XFILLER_11_483 VDD VSS sg13g2_decap_8
XFILLER_8_966 VDD VSS sg13g2_decap_8
XFILLER_23_91 VDD VSS sg13g2_decap_8
XFILLER_7_476 VDD VSS sg13g2_decap_8
XFILLER_48_1002 VDD VSS sg13g2_decap_8
XFILLER_98_704 VDD VSS sg13g2_decap_8
XFILLER_99_84 VDD VSS sg13g2_decap_8
XFILLER_98_748 VDD VSS sg13g2_fill_2
XFILLER_112_525 VDD VSS sg13g2_decap_8
XFILLER_97_214 VDD VSS sg13g2_decap_8
X_2300_ _2300_/RESET_B VSS VDD _2300_/D _2300_/Q _2368_/CLK sg13g2_dfrbpq_1
X_2231_ _2231_/RESET_B VSS VDD _2231_/D _2231_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_3_693 VDD VSS sg13g2_decap_8
XFILLER_78_450 VDD VSS sg13g2_decap_4
XFILLER_78_461 VDD VSS sg13g2_decap_8
XFILLER_39_815 VDD VSS sg13g2_decap_8
X_2162_ _2162_/A _2162_/B _2350_/D VDD VSS sg13g2_nor2_1
XFILLER_66_623 VDD VSS sg13g2_decap_8
XFILLER_94_976 VDD VSS sg13g2_decap_8
XFILLER_81_615 VDD VSS sg13g2_decap_8
XFILLER_93_442 VDD VSS sg13g2_decap_8
XFILLER_54_829 VDD VSS sg13g2_decap_8
XFILLER_53_306 VDD VSS sg13g2_decap_4
XFILLER_38_369 VDD VSS sg13g2_decap_8
X_2093_ _2093_/A _2093_/B _2094_/B VDD VSS sg13g2_nor2_1
XFILLER_94_1011 VDD VSS sg13g2_decap_8
XFILLER_65_177 VDD VSS sg13g2_decap_8
XFILLER_0_1015 VDD VSS sg13g2_decap_8
XFILLER_81_659 VDD VSS sg13g2_fill_1
XFILLER_34_553 VDD VSS sg13g2_decap_8
XFILLER_0_84 VDD VSS sg13g2_decap_8
XFILLER_94_1055 VDD VSS sg13g2_decap_4
XFILLER_61_361 VDD VSS sg13g2_fill_2
XFILLER_21_203 VDD VSS sg13g2_decap_8
X_1946_ _1946_/B _1946_/A _1984_/B VDD VSS sg13g2_xor2_1
XFILLER_30_770 VDD VSS sg13g2_decap_8
XFILLER_107_319 VDD VSS sg13g2_decap_4
X_1877_ _1877_/B _1877_/A _1879_/A VDD VSS sg13g2_xor2_1
XFILLER_31_1050 VDD VSS sg13g2_decap_8
XFILLER_103_503 VDD VSS sg13g2_decap_8
XFILLER_85_921 VDD VSS sg13g2_decap_4
XFILLER_88_269 VDD VSS sg13g2_decap_8
XFILLER_28_14 VDD VSS sg13g2_decap_8
XFILLER_85_943 VDD VSS sg13g2_decap_8
XFILLER_97_792 VDD VSS sg13g2_decap_4
XFILLER_96_280 VDD VSS sg13g2_decap_8
XFILLER_69_494 VDD VSS sg13g2_decap_8
XFILLER_29_336 VDD VSS sg13g2_decap_8
XFILLER_85_987 VDD VSS sg13g2_decap_4
XFILLER_57_667 VDD VSS sg13g2_decap_8
XFILLER_72_648 VDD VSS sg13g2_decap_8
XFILLER_72_615 VDD VSS sg13g2_decap_8
XFILLER_84_475 VDD VSS sg13g2_fill_1
XFILLER_38_870 VDD VSS sg13g2_decap_8
XFILLER_56_166 VDD VSS sg13g2_decap_8
XFILLER_44_35 VDD VSS sg13g2_decap_8
XFILLER_71_169 VDD VSS sg13g2_decap_8
XFILLER_53_873 VDD VSS sg13g2_decap_8
XFILLER_25_553 VDD VSS sg13g2_decap_8
XFILLER_12_203 VDD VSS sg13g2_decap_8
XFILLER_80_692 VDD VSS sg13g2_decap_4
XFILLER_40_512 VDD VSS sg13g2_decap_8
XFILLER_100_63 VDD VSS sg13g2_decap_8
XFILLER_40_578 VDD VSS sg13g2_decap_8
XFILLER_21_770 VDD VSS sg13g2_decap_8
XFILLER_60_45 VDD VSS sg13g2_decap_8
XFILLER_20_280 VDD VSS sg13g2_decap_8
XFILLER_5_903 VDD VSS sg13g2_decap_8
XFILLER_4_413 VDD VSS sg13g2_decap_8
XFILLER_107_842 VDD VSS sg13g2_decap_8
XFILLER_69_21 VDD VSS sg13g2_decap_8
XFILLER_79_203 VDD VSS sg13g2_decap_8
XFILLER_95_707 VDD VSS sg13g2_decap_8
XFILLER_0_630 VDD VSS sg13g2_decap_8
XFILLER_94_217 VDD VSS sg13g2_fill_1
XFILLER_88_781 VDD VSS sg13g2_decap_8
XFILLER_85_42 VDD VSS sg13g2_decap_8
XFILLER_48_645 VDD VSS sg13g2_decap_8
XFILLER_78_1028 VDD VSS sg13g2_decap_8
XFILLER_76_998 VDD VSS sg13g2_decap_4
XFILLER_75_486 VDD VSS sg13g2_decap_8
XFILLER_47_177 VDD VSS sg13g2_decap_8
XFILLER_44_851 VDD VSS sg13g2_decap_8
XFILLER_18_91 VDD VSS sg13g2_decap_8
XFILLER_62_169 VDD VSS sg13g2_decap_8
XFILLER_16_553 VDD VSS sg13g2_decap_8
XFILLER_43_350 VDD VSS sg13g2_decap_8
XFILLER_93_7 VDD VSS sg13g2_decap_8
X_1800_ _1811_/A _1800_/C _1800_/Y VDD VSS _1812_/B sg13g2_nand3b_1
XFILLER_54_1050 VDD VSS sg13g2_decap_8
XFILLER_31_567 VDD VSS sg13g2_decap_8
XFILLER_15_1001 VDD VSS sg13g2_decap_8
XFILLER_12_770 VDD VSS sg13g2_decap_8
X_1731_ _2235_/Q _2227_/Q _1926_/A VDD VSS sg13g2_nor2b_1
XFILLER_11_280 VDD VSS sg13g2_decap_8
XFILLER_8_763 VDD VSS sg13g2_decap_8
XFILLER_102_1059 VDD VSS sg13g2_fill_2
XFILLER_102_1048 VDD VSS sg13g2_decap_8
X_1662_ _2310_/Q _2333_/Q _2325_/Q _2348_/Q _2340_/Q _2311_/Q _1662_/X VDD VSS sg13g2_mux4_1
XFILLER_7_273 VDD VSS sg13g2_decap_8
X_2209__122 VDD VSS _2209_/RESET_B sg13g2_tiehi
XFILLER_4_980 VDD VSS sg13g2_decap_8
X_1593_ _1595_/A _1593_/B _1594_/B _2288_/D VDD VSS sg13g2_nor3_1
XFILLER_86_707 VDD VSS sg13g2_decap_4
XFILLER_112_322 VDD VSS sg13g2_decap_8
XFILLER_3_490 VDD VSS sg13g2_decap_8
XFILLER_98_567 VDD VSS sg13g2_decap_8
XFILLER_100_517 VDD VSS sg13g2_decap_8
XFILLER_85_217 VDD VSS sg13g2_decap_8
XFILLER_67_910 VDD VSS sg13g2_decap_8
XFILLER_112_399 VDD VSS sg13g2_decap_8
X_2214_ _2214_/RESET_B VSS VDD _2214_/D _2214_/Q clkload7/A sg13g2_dfrbpq_1
XFILLER_67_921 VDD VSS sg13g2_fill_1
XFILLER_67_932 VDD VSS sg13g2_fill_1
XFILLER_61_1054 VDD VSS sg13g2_decap_8
XFILLER_39_612 VDD VSS sg13g2_decap_8
X_2145_ VDD VSS _2124_/B _2120_/A _2144_/X hold312/X _2147_/A _2124_/Y sg13g2_a221oi_1
XFILLER_66_442 VDD VSS sg13g2_decap_8
XFILLER_15_0 VDD VSS sg13g2_decap_8
XFILLER_38_133 VDD VSS sg13g2_decap_8
XFILLER_82_935 VDD VSS sg13g2_decap_8
XFILLER_81_412 VDD VSS sg13g2_decap_8
XFILLER_39_689 VDD VSS sg13g2_decap_8
X_2076_ _2076_/Y _2082_/B _2076_/B VDD VSS sg13g2_nand2_1
XFILLER_35_840 VDD VSS sg13g2_decap_8
XFILLER_81_489 VDD VSS sg13g2_decap_8
XFILLER_34_350 VDD VSS sg13g2_decap_8
XFILLER_50_887 VDD VSS sg13g2_decap_8
XFILLER_22_567 VDD VSS sg13g2_decap_8
XFILLER_14_49 VDD VSS sg13g2_decap_8
XFILLER_10_707 VDD VSS sg13g2_decap_8
X_1929_ _1931_/A _1929_/A _1929_/B VDD VSS sg13g2_xnor2_1
XFILLER_107_105 VDD VSS sg13g2_decap_8
Xfanout1 _2162_/B _2156_/A VDD VSS sg13g2_buf_1
XFILLER_89_501 VDD VSS sg13g2_decap_8
XFILLER_2_917 VDD VSS sg13g2_decap_8
XFILLER_104_834 VDD VSS sg13g2_decap_4
XFILLER_1_427 VDD VSS sg13g2_decap_8
XFILLER_103_355 VDD VSS sg13g2_decap_8
XFILLER_39_35 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[4\].out_data_pad out_data_PADs[4] bondpad_70x70
XFILLER_58_943 VDD VSS sg13g2_decap_8
XFILLER_85_751 VDD VSS sg13g2_fill_1
XFILLER_58_987 VDD VSS sg13g2_decap_8
XFILLER_57_453 VDD VSS sg13g2_decap_8
XFILLER_29_133 VDD VSS sg13g2_decap_8
XFILLER_85_784 VDD VSS sg13g2_decap_8
XFILLER_45_637 VDD VSS sg13g2_decap_4
XFILLER_57_464 VDD VSS sg13g2_fill_2
XFILLER_26_840 VDD VSS sg13g2_decap_8
XFILLER_55_56 VDD VSS sg13g2_decap_8
XFILLER_25_350 VDD VSS sg13g2_decap_8
XFILLER_38_1045 VDD VSS sg13g2_decap_8
XFILLER_41_832 VDD VSS sg13g2_decap_8
XFILLER_111_84 VDD VSS sg13g2_decap_8
XFILLER_13_567 VDD VSS sg13g2_decap_8
XFILLER_40_342 VDD VSS sg13g2_decap_8
XFILLER_71_88 VDD VSS sg13g2_decap_4
XFILLER_5_700 VDD VSS sg13g2_decap_8
XFILLER_4_210 VDD VSS sg13g2_decap_8
XFILLER_20_70 VDD VSS sg13g2_decap_8
XFILLER_5_777 VDD VSS sg13g2_decap_8
XFILLER_106_182 VDD VSS sg13g2_decap_8
XFILLER_4_287 VDD VSS sg13g2_decap_8
XFILLER_95_515 VDD VSS sg13g2_decap_8
XFILLER_45_1038 VDD VSS sg13g2_decap_8
XFILLER_68_729 VDD VSS sg13g2_decap_4
XFILLER_110_837 VDD VSS sg13g2_decap_8
XFILLER_96_63 VDD VSS sg13g2_decap_8
XFILLER_1_994 VDD VSS sg13g2_decap_8
XFILLER_76_762 VDD VSS sg13g2_decap_8
XFILLER_75_250 VDD VSS sg13g2_decap_8
XFILLER_36_637 VDD VSS sg13g2_decap_8
XFILLER_63_401 VDD VSS sg13g2_decap_8
XFILLER_17_840 VDD VSS sg13g2_decap_8
XFILLER_35_147 VDD VSS sg13g2_decap_8
XFILLER_91_787 VDD VSS sg13g2_decap_8
XFILLER_90_242 VDD VSS sg13g2_decap_8
XFILLER_63_489 VDD VSS sg13g2_decap_8
XFILLER_16_350 VDD VSS sg13g2_decap_8
XFILLER_50_106 VDD VSS sg13g2_decap_8
XFILLER_91_1014 VDD VSS sg13g2_decap_8
XFILLER_72_990 VDD VSS sg13g2_decap_8
XFILLER_32_854 VDD VSS sg13g2_decap_8
XFILLER_31_364 VDD VSS sg13g2_decap_8
X_1714_ _1719_/B _1714_/A _1723_/B VDD VSS sg13g2_xnor2_1
XFILLER_8_560 VDD VSS sg13g2_decap_8
XFILLER_105_609 VDD VSS sg13g2_decap_8
XFILLER_99_810 VDD VSS sg13g2_fill_1
XFILLER_104_119 VDD VSS sg13g2_decap_8
X_1645_ _2298_/D _1645_/B _2307_/D VDD VSS sg13g2_nand2b_1
XFILLER_99_843 VDD VSS sg13g2_decap_8
X_1576_ _1576_/A _1576_/B _2281_/D VDD VSS sg13g2_nor2_1
XFILLER_98_353 VDD VSS sg13g2_decap_8
XFILLER_100_314 VDD VSS sg13g2_decap_8
XFILLER_98_397 VDD VSS sg13g2_decap_8
XFILLER_112_196 VDD VSS sg13g2_decap_8
XFILLER_67_762 VDD VSS sg13g2_decap_8
XFILLER_67_740 VDD VSS sg13g2_fill_2
XFILLER_55_902 VDD VSS sg13g2_decap_8
XFILLER_6_1043 VDD VSS sg13g2_decap_8
XFILLER_39_464 VDD VSS sg13g2_decap_8
X_2128_ _2124_/A _2198_/Q _2190_/Q _2182_/Q _2174_/Q _2144_/S1 _2128_/X VDD VSS sg13g2_mux4_1
XFILLER_27_637 VDD VSS sg13g2_decap_8
XFILLER_66_294 VDD VSS sg13g2_decap_8
X_2257__237 VDD VSS _2257_/RESET_B sg13g2_tiehi
XFILLER_70_927 VDD VSS sg13g2_decap_8
XFILLER_82_765 VDD VSS sg13g2_fill_2
X_2059_ _2059_/Y _2074_/A _2083_/A VDD VSS sg13g2_nand2_1
XFILLER_81_242 VDD VSS sg13g2_decap_8
XFILLER_54_467 VDD VSS sg13g2_decap_8
XFILLER_26_147 VDD VSS sg13g2_decap_8
XFILLER_23_854 VDD VSS sg13g2_decap_8
XFILLER_10_504 VDD VSS sg13g2_decap_8
XFILLER_41_14 VDD VSS sg13g2_decap_8
XFILLER_22_364 VDD VSS sg13g2_decap_8
XFILLER_109_959 VDD VSS sg13g2_decap_8
XFILLER_108_436 VDD VSS sg13g2_decap_8
XFILLER_2_714 VDD VSS sg13g2_decap_8
Xhold560 _1725_/Y VDD VSS _2320_/D sg13g2_dlygate4sd3_1
XFILLER_1_224 VDD VSS sg13g2_decap_8
XFILLER_104_675 VDD VSS sg13g2_decap_8
XFILLER_89_342 VDD VSS sg13g2_decap_8
XFILLER_77_537 VDD VSS sg13g2_decap_8
XFILLER_49_239 VDD VSS sg13g2_decap_8
XFILLER_103_196 VDD VSS sg13g2_decap_8
XFILLER_106_84 VDD VSS sg13g2_decap_8
XFILLER_58_795 VDD VSS sg13g2_decap_8
XFILLER_66_77 VDD VSS sg13g2_decap_8
XFILLER_46_968 VDD VSS sg13g2_decap_8
XFILLER_57_283 VDD VSS sg13g2_decap_8
XFILLER_18_637 VDD VSS sg13g2_decap_8
XFILLER_82_21 VDD VSS sg13g2_decap_8
XFILLER_17_147 VDD VSS sg13g2_decap_8
XFILLER_54_990 VDD VSS sg13g2_decap_8
XFILLER_82_98 VDD VSS sg13g2_decap_8
XFILLER_14_854 VDD VSS sg13g2_decap_8
XFILLER_13_364 VDD VSS sg13g2_decap_8
XFILLER_15_70 VDD VSS sg13g2_decap_8
XFILLER_40_161 VDD VSS sg13g2_decap_8
XFILLER_51_1031 VDD VSS sg13g2_decap_8
XFILLER_9_357 VDD VSS sg13g2_decap_8
XFILLER_12_1015 VDD VSS sg13g2_decap_8
XFILLER_5_574 VDD VSS sg13g2_decap_8
XFILLER_31_91 VDD VSS sg13g2_decap_8
XFILLER_56_7 VDD VSS sg13g2_decap_8
X_1430_ _1431_/A _1429_/Y hold469/X _1429_/B _1364_/A VDD VSS sg13g2_a22oi_1
X_1361_ VDD _2209_/D _1361_/A VSS sg13g2_inv_1
XFILLER_110_634 VDD VSS sg13g2_decap_8
XFILLER_96_857 VDD VSS sg13g2_decap_8
XFILLER_68_537 VDD VSS sg13g2_decap_8
XFILLER_68_515 VDD VSS sg13g2_decap_4
X_1292_ _1292_/Y _1342_/B1 hold357/X _1342_/A2 _2340_/Q VDD VSS sg13g2_a22oi_1
XFILLER_1_791 VDD VSS sg13g2_decap_8
XFILLER_83_529 VDD VSS sg13g2_decap_8
XFILLER_83_518 VDD VSS sg13g2_fill_2
XFILLER_37_924 VDD VSS sg13g2_decap_8
XFILLER_49_762 VDD VSS sg13g2_decap_8
XFILLER_64_732 VDD VSS sg13g2_decap_8
XFILLER_36_434 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_91_584 VDD VSS sg13g2_decap_8
XFILLER_63_297 VDD VSS sg13g2_decap_8
XFILLER_51_415 VDD VSS sg13g2_decap_8
XFILLER_108_1032 VDD VSS sg13g2_decap_8
XFILLER_32_651 VDD VSS sg13g2_decap_8
XFILLER_31_161 VDD VSS sg13g2_decap_8
XFILLER_82_0 VDD VSS sg13g2_decap_8
XFILLER_20_868 VDD VSS sg13g2_decap_8
XFILLER_11_28 VDD VSS sg13g2_decap_8
XFILLER_105_428 VDD VSS sg13g2_decap_8
X_1628_ _1633_/B _1628_/A _1637_/B VDD VSS sg13g2_xnor2_1
XFILLER_99_673 VDD VSS sg13g2_decap_8
XFILLER_67_1060 VDD VSS sg13g2_fill_1
XFILLER_28_1022 VDD VSS sg13g2_decap_8
XFILLER_59_504 VDD VSS sg13g2_decap_8
XFILLER_101_601 VDD VSS sg13g2_decap_8
XFILLER_98_183 VDD VSS sg13g2_decap_8
X_1559_ _1558_/Y VDD _1559_/Y VSS _1573_/A1 _2207_/Q sg13g2_o21ai_1
XFILLER_87_857 VDD VSS sg13g2_decap_8
XFILLER_86_356 VDD VSS sg13g2_decap_8
XFILLER_100_133 VDD VSS sg13g2_decap_8
XFILLER_101_678 VDD VSS sg13g2_decap_8
XFILLER_100_166 VDD VSS sg13g2_fill_1
XFILLER_74_518 VDD VSS sg13g2_decap_8
XFILLER_74_507 VDD VSS sg13g2_decap_8
XFILLER_28_924 VDD VSS sg13g2_decap_8
XFILLER_67_581 VDD VSS sg13g2_decap_8
XFILLER_54_220 VDD VSS sg13g2_decap_8
XFILLER_36_14 VDD VSS sg13g2_decap_8
XFILLER_27_434 VDD VSS sg13g2_decap_8
XFILLER_82_562 VDD VSS sg13g2_decap_8
XFILLER_55_776 VDD VSS sg13g2_fill_2
XFILLER_43_905 VDD VSS sg13g2_decap_8
XFILLER_70_724 VDD VSS sg13g2_decap_8
XFILLER_54_275 VDD VSS sg13g2_fill_1
XFILLER_42_426 VDD VSS sg13g2_decap_8
XFILLER_74_1031 VDD VSS sg13g2_decap_8
XFILLER_23_651 VDD VSS sg13g2_decap_8
XFILLER_51_982 VDD VSS sg13g2_decap_8
XFILLER_35_1015 VDD VSS sg13g2_decap_8
XFILLER_10_301 VDD VSS sg13g2_decap_8
XFILLER_22_161 VDD VSS sg13g2_decap_8
X_2311__286 VDD VSS _2311_/RESET_B sg13g2_tiehi
XFILLER_11_868 VDD VSS sg13g2_decap_8
XFILLER_109_756 VDD VSS sg13g2_decap_8
XFILLER_108_222 VDD VSS sg13g2_decap_8
XFILLER_10_378 VDD VSS sg13g2_decap_8
XFILLER_2_511 VDD VSS sg13g2_decap_8
XFILLER_105_973 VDD VSS sg13g2_decap_8
XFILLER_78_813 VDD VSS sg13g2_decap_8
XFILLER_77_21 VDD VSS sg13g2_decap_8
Xhold390 _1316_/Y VDD VSS _1317_/A sg13g2_dlygate4sd3_1
XFILLER_104_472 VDD VSS sg13g2_decap_4
XFILLER_77_301 VDD VSS sg13g2_decap_8
XFILLER_89_161 VDD VSS sg13g2_decap_8
XFILLER_42_1008 VDD VSS sg13g2_decap_8
XFILLER_2_588 VDD VSS sg13g2_decap_8
XFILLER_77_98 VDD VSS sg13g2_decap_8
XFILLER_58_570 VDD VSS sg13g2_decap_8
XFILLER_46_710 VDD VSS sg13g2_decap_4
XFILLER_65_529 VDD VSS sg13g2_decap_8
XFILLER_19_924 VDD VSS sg13g2_decap_8
XFILLER_92_326 VDD VSS sg13g2_decap_8
XFILLER_93_42 VDD VSS sg13g2_decap_8
XFILLER_18_434 VDD VSS sg13g2_decap_8
XFILLER_46_754 VDD VSS sg13g2_decap_8
XFILLER_34_938 VDD VSS sg13g2_decap_8
XFILLER_61_735 VDD VSS sg13g2_fill_2
XFILLER_61_779 VDD VSS sg13g2_decap_4
XFILLER_60_256 VDD VSS sg13g2_decap_8
XFILLER_26_91 VDD VSS sg13g2_decap_8
XFILLER_33_448 VDD VSS sg13g2_decap_8
XFILLER_14_651 VDD VSS sg13g2_decap_8
XFILLER_13_161 VDD VSS sg13g2_decap_8
X_2171__198 VDD VSS _2171_/RESET_B sg13g2_tiehi
XFILLER_9_154 VDD VSS sg13g2_decap_8
XFILLER_6_861 VDD VSS sg13g2_decap_8
XFILLER_5_371 VDD VSS sg13g2_decap_8
XFILLER_87_109 VDD VSS sg13g2_decap_8
XFILLER_111_910 VDD VSS sg13g2_decap_8
X_1413_ _1412_/Y VDD _2227_/D VSS _1364_/Y _1410_/Y sg13g2_o21ai_1
XFILLER_68_312 VDD VSS sg13g2_decap_8
XFILLER_96_665 VDD VSS sg13g2_decap_8
XFILLER_69_868 VDD VSS sg13g2_decap_8
XFILLER_110_431 VDD VSS sg13g2_decap_8
X_1344_ _1344_/Y _1344_/B1 hold353/X _1344_/A2 _2335_/Q VDD VSS sg13g2_a22oi_1
XFILLER_111_987 VDD VSS sg13g2_decap_8
X_1275_ VDD _2167_/D _1275_/A VSS sg13g2_inv_1
XFILLER_95_175 VDD VSS sg13g2_decap_8
XFILLER_3_84 VDD VSS sg13g2_decap_8
XFILLER_37_721 VDD VSS sg13g2_decap_8
XFILLER_58_1015 VDD VSS sg13g2_decap_4
XFILLER_3_1057 VDD VSS sg13g2_decap_4
XFILLER_36_231 VDD VSS sg13g2_decap_8
XFILLER_25_938 VDD VSS sg13g2_decap_8
XFILLER_37_798 VDD VSS sg13g2_decap_8
XFILLER_58_1059 VDD VSS sg13g2_fill_2
XFILLER_52_779 VDD VSS sg13g2_decap_4
XFILLER_24_448 VDD VSS sg13g2_decap_8
XFILLER_51_223 VDD VSS sg13g2_decap_8
XFILLER_20_665 VDD VSS sg13g2_decap_8
XFILLER_22_49 VDD VSS sg13g2_decap_8
XFILLER_3_308 VDD VSS sg13g2_decap_8
XFILLER_106_748 VDD VSS sg13g2_decap_8
XFILLER_65_1008 VDD VSS sg13g2_decap_8
XFILLER_59_312 VDD VSS sg13g2_fill_2
XFILLER_59_334 VDD VSS sg13g2_decap_8
XFILLER_75_827 VDD VSS sg13g2_decap_8
XFILLER_86_164 VDD VSS sg13g2_decap_8
XFILLER_47_35 VDD VSS sg13g2_decap_8
XFILLER_101_486 VDD VSS sg13g2_decap_4
XFILLER_68_890 VDD VSS sg13g2_decap_8
XFILLER_28_721 VDD VSS sg13g2_decap_8
XFILLER_83_871 VDD VSS sg13g2_decap_8
XFILLER_74_359 VDD VSS sg13g2_decap_8
XFILLER_43_702 VDD VSS sg13g2_decap_8
XFILLER_55_540 VDD VSS sg13g2_fill_2
XFILLER_27_231 VDD VSS sg13g2_decap_8
XFILLER_103_63 VDD VSS sg13g2_decap_8
XFILLER_55_595 VDD VSS sg13g2_fill_2
XFILLER_28_798 VDD VSS sg13g2_decap_8
XFILLER_16_938 VDD VSS sg13g2_decap_8
XFILLER_42_212 VDD VSS sg13g2_decap_8
XFILLER_15_448 VDD VSS sg13g2_decap_8
XFILLER_63_56 VDD VSS sg13g2_decap_8
XFILLER_42_245 VDD VSS sg13g2_decap_8
XFILLER_43_779 VDD VSS sg13g2_decap_8
XFILLER_70_598 VDD VSS sg13g2_decap_8
XFILLER_11_665 VDD VSS sg13g2_decap_8
XFILLER_10_175 VDD VSS sg13g2_decap_8
XFILLER_7_658 VDD VSS sg13g2_decap_8
XFILLER_109_553 VDD VSS sg13g2_decap_8
XFILLER_6_168 VDD VSS sg13g2_decap_8
XFILLER_112_707 VDD VSS sg13g2_decap_8
XFILLER_97_407 VDD VSS sg13g2_decap_8
XFILLER_88_42 VDD VSS sg13g2_decap_8
XFILLER_105_770 VDD VSS sg13g2_decap_8
XFILLER_78_621 VDD VSS sg13g2_decap_8
XFILLER_111_217 VDD VSS sg13g2_decap_8
XFILLER_3_875 VDD VSS sg13g2_decap_8
XFILLER_104_280 VDD VSS sg13g2_decap_8
XFILLER_2_385 VDD VSS sg13g2_decap_8
XFILLER_66_838 VDD VSS sg13g2_decap_4
XFILLER_93_635 VDD VSS sg13g2_decap_8
XFILLER_77_175 VDD VSS sg13g2_decap_8
XFILLER_92_112 VDD VSS sg13g2_fill_1
XFILLER_19_7 VDD VSS sg13g2_decap_8
XFILLER_19_721 VDD VSS sg13g2_decap_8
XFILLER_93_679 VDD VSS sg13g2_decap_4
XFILLER_81_819 VDD VSS sg13g2_fill_2
XFILLER_81_808 VDD VSS sg13g2_decap_8
XFILLER_46_551 VDD VSS sg13g2_fill_1
XFILLER_18_231 VDD VSS sg13g2_decap_8
XFILLER_92_178 VDD VSS sg13g2_decap_8
XFILLER_34_735 VDD VSS sg13g2_decap_8
XFILLER_19_798 VDD VSS sg13g2_decap_8
X_2357__275 VDD VSS _2357_/RESET_B sg13g2_tiehi
XFILLER_61_543 VDD VSS sg13g2_decap_8
XFILLER_33_245 VDD VSS sg13g2_decap_8
X_1962_ _1962_/B _1962_/A _1982_/B VDD VSS sg13g2_xor2_1
XFILLER_18_1043 VDD VSS sg13g2_decap_8
X_1893_ _1892_/B _1892_/X _1954_/S _1960_/B VDD VSS sg13g2_mux2_1
XFILLER_30_952 VDD VSS sg13g2_decap_8
XFILLER_105_1057 VDD VSS sg13g2_decap_4
XFILLER_89_908 VDD VSS sg13g2_decap_8
XFILLER_45_0 VDD VSS sg13g2_decap_8
XFILLER_97_930 VDD VSS sg13g2_decap_8
XFILLER_69_621 VDD VSS sg13g2_decap_8
XFILLER_88_429 VDD VSS sg13g2_decap_8
XFILLER_84_613 VDD VSS sg13g2_decap_8
XFILLER_96_473 VDD VSS sg13g2_fill_2
XFILLER_96_462 VDD VSS sg13g2_decap_8
XFILLER_25_1036 VDD VSS sg13g2_decap_8
XFILLER_29_518 VDD VSS sg13g2_decap_8
XFILLER_111_784 VDD VSS sg13g2_decap_8
X_1327_ VDD _2193_/D _1327_/A VSS sg13g2_inv_1
XFILLER_83_112 VDD VSS sg13g2_decap_8
XFILLER_68_197 VDD VSS sg13g2_decap_8
XFILLER_56_326 VDD VSS sg13g2_decap_8
XFILLER_72_808 VDD VSS sg13g2_fill_2
XFILLER_110_294 VDD VSS sg13g2_decap_8
X_1258_ VSS VDD _1265_/B _1257_/Y _1258_/Y _1228_/A sg13g2_a21oi_1
X_2219__102 VDD VSS _2219_/RESET_B sg13g2_tiehi
X_1189_ VDD _1189_/Y _2298_/Q VSS sg13g2_inv_1
XFILLER_25_735 VDD VSS sg13g2_decap_8
XFILLER_17_49 VDD VSS sg13g2_decap_8
XFILLER_37_595 VDD VSS sg13g2_decap_8
XFILLER_64_381 VDD VSS sg13g2_decap_8
XFILLER_24_245 VDD VSS sg13g2_decap_8
XFILLER_52_576 VDD VSS sg13g2_decap_8
XFILLER_71_1012 VDD VSS sg13g2_decap_8
XFILLER_21_952 VDD VSS sg13g2_decap_8
XFILLER_32_1029 VDD VSS sg13g2_decap_8
XFILLER_20_462 VDD VSS sg13g2_decap_8
XFILLER_3_105 VDD VSS sg13g2_decap_8
Xout_data_pads\[1\].out_data_pad _2367_/Q IOVDD IOVSS out_data_PADs[1] VDD VSS sg13g2_IOPadOut30mA
XFILLER_0_812 VDD VSS sg13g2_decap_8
XFILLER_102_773 VDD VSS sg13g2_decap_8
XFILLER_75_602 VDD VSS sg13g2_decap_8
XFILLER_87_451 VDD VSS sg13g2_decap_8
XFILLER_87_462 VDD VSS sg13g2_fill_2
XFILLER_0_889 VDD VSS sg13g2_decap_8
XFILLER_59_131 VDD VSS sg13g2_fill_2
XFILLER_102_795 VDD VSS sg13g2_decap_8
XFILLER_101_283 VDD VSS sg13g2_decap_8
XFILLER_74_112 VDD VSS sg13g2_decap_8
XFILLER_75_679 VDD VSS sg13g2_decap_8
XFILLER_74_77 VDD VSS sg13g2_decap_8
XFILLER_56_871 VDD VSS sg13g2_decap_8
XFILLER_28_595 VDD VSS sg13g2_decap_8
XFILLER_55_392 VDD VSS sg13g2_decap_8
XFILLER_16_735 VDD VSS sg13g2_decap_8
XFILLER_43_521 VDD VSS sg13g2_decap_8
XFILLER_70_351 VDD VSS sg13g2_decap_8
X_2237__268 VDD VSS _2237_/RESET_B sg13g2_tiehi
XFILLER_90_21 VDD VSS sg13g2_decap_8
XFILLER_43_576 VDD VSS sg13g2_decap_8
XFILLER_15_245 VDD VSS sg13g2_decap_8
XFILLER_31_749 VDD VSS sg13g2_decap_8
XFILLER_12_952 VDD VSS sg13g2_decap_8
XFILLER_30_259 VDD VSS sg13g2_decap_8
XFILLER_90_98 VDD VSS sg13g2_decap_8
XFILLER_11_462 VDD VSS sg13g2_decap_8
XFILLER_8_945 VDD VSS sg13g2_decap_8
XFILLER_23_70 VDD VSS sg13g2_decap_8
XFILLER_7_455 VDD VSS sg13g2_decap_8
XFILLER_99_63 VDD VSS sg13g2_decap_8
XFILLER_112_504 VDD VSS sg13g2_decap_8
XFILLER_48_1058 VDD VSS sg13g2_fill_2
XFILLER_3_672 VDD VSS sg13g2_decap_8
X_2230_ _2230__80/L_HI VSS VDD _2230_/D _2230_/Q clkload6/A sg13g2_dfrbpq_1
XFILLER_2_182 VDD VSS sg13g2_decap_8
XFILLER_94_955 VDD VSS sg13g2_decap_8
XFILLER_93_421 VDD VSS sg13g2_decap_8
X_2161_ _2162_/A _2162_/B _2349_/D VDD VSS sg13g2_nor2_1
XFILLER_65_112 VDD VSS sg13g2_fill_2
XFILLER_65_101 VDD VSS sg13g2_decap_8
XFILLER_54_808 VDD VSS sg13g2_decap_8
XFILLER_65_156 VDD VSS sg13g2_decap_8
XFILLER_38_348 VDD VSS sg13g2_decap_8
X_2092_ _2092_/A _1252_/Y _2102_/B VDD VSS sg13g2_nor2b_1
XFILLER_111_1050 VDD VSS sg13g2_decap_8
XFILLER_93_498 VDD VSS sg13g2_decap_8
XFILLER_94_1034 VDD VSS sg13g2_decap_8
XFILLER_0_63 VDD VSS sg13g2_decap_8
XFILLER_19_595 VDD VSS sg13g2_decap_8
XFILLER_34_532 VDD VSS sg13g2_decap_8
XFILLER_62_885 VDD VSS sg13g2_decap_8
XFILLER_22_749 VDD VSS sg13g2_decap_8
X_1945_ _1946_/A _1946_/B _1945_/X VDD VSS sg13g2_and2_1
XFILLER_21_259 VDD VSS sg13g2_decap_8
X_1876_ _1876_/A _1876_/B _1971_/A VDD VSS sg13g2_and2_1
XFILLER_1_609 VDD VSS sg13g2_decap_8
XFILLER_103_537 VDD VSS sg13g2_decap_8
XFILLER_88_248 VDD VSS sg13g2_decap_8
XFILLER_0_119 VDD VSS sg13g2_decap_8
XFILLER_97_771 VDD VSS sg13g2_decap_8
XFILLER_111_581 VDD VSS sg13g2_decap_8
XFILLER_69_473 VDD VSS sg13g2_decap_8
XFILLER_57_646 VDD VSS sg13g2_decap_8
X_2359_ _2359_/RESET_B VSS VDD _2359_/D _2359_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_29_315 VDD VSS sg13g2_decap_8
XFILLER_56_145 VDD VSS sg13g2_decap_8
XFILLER_72_627 VDD VSS sg13g2_decap_8
XFILLER_44_329 VDD VSS sg13g2_decap_8
XFILLER_71_148 VDD VSS sg13g2_decap_8
XFILLER_53_852 VDD VSS sg13g2_decap_8
XFILLER_44_14 VDD VSS sg13g2_decap_8
XFILLER_25_532 VDD VSS sg13g2_decap_8
XFILLER_37_392 VDD VSS sg13g2_decap_8
XFILLER_80_671 VDD VSS sg13g2_decap_8
XFILLER_13_749 VDD VSS sg13g2_decap_8
XFILLER_40_535 VDD VSS sg13g2_fill_2
XFILLER_100_42 VDD VSS sg13g2_decap_8
XFILLER_40_557 VDD VSS sg13g2_decap_8
XFILLER_12_259 VDD VSS sg13g2_decap_8
XFILLER_107_821 VDD VSS sg13g2_decap_8
XFILLER_5_959 VDD VSS sg13g2_decap_8
XFILLER_107_898 VDD VSS sg13g2_decap_8
XFILLER_109_84 VDD VSS sg13g2_decap_8
XFILLER_4_469 VDD VSS sg13g2_decap_8
XFILLER_106_386 VDD VSS sg13g2_decap_8
XFILLER_69_99 VDD VSS sg13g2_decap_8
XFILLER_76_900 VDD VSS sg13g2_decap_8
XFILLER_102_581 VDD VSS sg13g2_decap_8
XFILLER_85_21 VDD VSS sg13g2_decap_8
XFILLER_48_624 VDD VSS sg13g2_decap_8
XFILLER_0_686 VDD VSS sg13g2_decap_8
XFILLER_76_977 VDD VSS sg13g2_decap_8
XFILLER_75_432 VDD VSS sg13g2_fill_1
XFILLER_36_819 VDD VSS sg13g2_decap_8
XFILLER_91_947 VDD VSS sg13g2_decap_8
XFILLER_75_465 VDD VSS sg13g2_decap_8
XFILLER_85_98 VDD VSS sg13g2_decap_8
XFILLER_29_882 VDD VSS sg13g2_decap_8
XFILLER_18_70 VDD VSS sg13g2_decap_8
XFILLER_35_329 VDD VSS sg13g2_decap_8
XFILLER_47_167 VDD VSS sg13g2_fill_1
XFILLER_90_424 VDD VSS sg13g2_decap_4
XFILLER_63_649 VDD VSS sg13g2_decap_8
XFILLER_16_532 VDD VSS sg13g2_decap_8
XFILLER_62_148 VDD VSS sg13g2_decap_8
XFILLER_28_392 VDD VSS sg13g2_decap_8
XFILLER_71_682 VDD VSS sg13g2_fill_2
Xin_valid_pad IOVDD IOVSS _1365_/B in_valid_PAD VDD VSS sg13g2_IOPadIn
XFILLER_31_546 VDD VSS sg13g2_decap_8
XFILLER_34_91 VDD VSS sg13g2_decap_8
XFILLER_86_7 VDD VSS sg13g2_decap_8
XFILLER_102_1027 VDD VSS sg13g2_decap_8
X_1730_ _1730_/Y _2236_/Q _2228_/Q VDD VSS sg13g2_nand2b_1
XFILLER_8_742 VDD VSS sg13g2_decap_8
XFILLER_15_1057 VDD VSS sg13g2_decap_4
X_1661_ _1670_/A _1661_/B _2303_/D VDD VSS sg13g2_nor2_1
XFILLER_7_252 VDD VSS sg13g2_decap_8
XFILLER_112_301 VDD VSS sg13g2_decap_8
X_1592_ _1592_/A _1592_/B _1594_/B VDD VSS sg13g2_and2_1
XIO_FILL_IO_EAST_6_2 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_98_546 VDD VSS sg13g2_decap_8
XFILLER_79_771 VDD VSS sg13g2_decap_8
XFILLER_112_378 VDD VSS sg13g2_decap_8
X_2213_ _2213_/RESET_B VSS VDD _2213_/D _2213_/Q _2245_/CLK sg13g2_dfrbpq_1
XFILLER_61_1033 VDD VSS sg13g2_decap_8
XFILLER_38_112 VDD VSS sg13g2_decap_8
X_2144_ _2144_/S0 _2202_/Q _2194_/Q _2186_/Q _2178_/Q _2144_/S1 _2144_/X VDD VSS sg13g2_mux4_1
XFILLER_39_668 VDD VSS sg13g2_decap_8
XFILLER_27_819 VDD VSS sg13g2_decap_8
XFILLER_82_914 VDD VSS sg13g2_decap_8
XFILLER_67_999 VDD VSS sg13g2_decap_8
XFILLER_53_104 VDD VSS sg13g2_decap_8
XFILLER_26_329 VDD VSS sg13g2_decap_8
X_2075_ _2076_/B _2075_/B _2004_/B VDD VSS sg13g2_nand2b_1
XFILLER_66_498 VDD VSS sg13g2_decap_8
XFILLER_19_392 VDD VSS sg13g2_decap_8
XFILLER_38_189 VDD VSS sg13g2_decap_8
XFILLER_81_468 VDD VSS sg13g2_decap_8
XFILLER_90_980 VDD VSS sg13g2_decap_8
XFILLER_62_693 VDD VSS sg13g2_decap_8
XFILLER_50_844 VDD VSS sg13g2_fill_1
XFILLER_50_833 VDD VSS sg13g2_decap_8
XFILLER_35_896 VDD VSS sg13g2_decap_8
XFILLER_22_546 VDD VSS sg13g2_decap_8
XFILLER_61_192 VDD VSS sg13g2_decap_8
XFILLER_14_28 VDD VSS sg13g2_decap_8
X_1928_ _1933_/A _1928_/A _1928_/B VDD VSS sg13g2_xnor2_1
X_1859_ _1934_/B _2003_/A _1907_/A VDD VSS sg13g2_and2_1
Xfanout2 _2160_/B _2162_/B VDD VSS sg13g2_buf_1
XFILLER_30_49 VDD VSS sg13g2_decap_8
XFILLER_104_813 VDD VSS sg13g2_decap_8
XFILLER_1_406 VDD VSS sg13g2_decap_8
XFILLER_103_334 VDD VSS sg13g2_decap_8
XFILLER_39_14 VDD VSS sg13g2_decap_8
XFILLER_76_207 VDD VSS sg13g2_fill_1
XFILLER_58_922 VDD VSS sg13g2_decap_8
XFILLER_29_112 VDD VSS sg13g2_decap_8
XFILLER_85_763 VDD VSS sg13g2_decap_8
XFILLER_69_281 VDD VSS sg13g2_decap_8
XFILLER_57_432 VDD VSS sg13g2_decap_8
XFILLER_18_819 VDD VSS sg13g2_decap_8
XFILLER_55_35 VDD VSS sg13g2_decap_8
XFILLER_17_329 VDD VSS sg13g2_decap_8
XFILLER_29_189 VDD VSS sg13g2_decap_8
XFILLER_60_619 VDD VSS sg13g2_decap_4
XFILLER_44_148 VDD VSS sg13g2_decap_8
XFILLER_81_991 VDD VSS sg13g2_fill_1
XFILLER_111_63 VDD VSS sg13g2_decap_8
XFILLER_38_1024 VDD VSS sg13g2_decap_8
XFILLER_41_811 VDD VSS sg13g2_decap_8
XFILLER_26_896 VDD VSS sg13g2_decap_8
XFILLER_71_56 VDD VSS sg13g2_decap_8
XFILLER_13_546 VDD VSS sg13g2_decap_8
XFILLER_40_321 VDD VSS sg13g2_decap_8
XFILLER_52_181 VDD VSS sg13g2_decap_8
XFILLER_41_888 VDD VSS sg13g2_decap_8
XFILLER_9_539 VDD VSS sg13g2_decap_8
XFILLER_40_398 VDD VSS sg13g2_decap_8
XFILLER_112_0 VDD VSS sg13g2_decap_8
XFILLER_5_756 VDD VSS sg13g2_decap_8
XFILLER_4_266 VDD VSS sg13g2_decap_8
XFILLER_84_1044 VDD VSS sg13g2_decap_8
XFILLER_107_695 VDD VSS sg13g2_decap_8
XFILLER_106_161 VDD VSS sg13g2_decap_8
XFILLER_45_1017 VDD VSS sg13g2_decap_8
XFILLER_110_816 VDD VSS sg13g2_decap_8
XFILLER_96_42 VDD VSS sg13g2_decap_8
XFILLER_68_708 VDD VSS sg13g2_decap_8
XFILLER_49_911 VDD VSS sg13g2_decap_8
XFILLER_1_973 VDD VSS sg13g2_decap_8
XFILLER_76_741 VDD VSS sg13g2_decap_8
XFILLER_0_483 VDD VSS sg13g2_decap_8
XFILLER_49_988 VDD VSS sg13g2_decap_8
XFILLER_36_616 VDD VSS sg13g2_decap_8
XFILLER_29_91 VDD VSS sg13g2_decap_8
XFILLER_64_958 VDD VSS sg13g2_decap_8
XFILLER_21_1050 VDD VSS sg13g2_decap_8
XFILLER_35_126 VDD VSS sg13g2_decap_8
XFILLER_91_766 VDD VSS sg13g2_decap_8
XFILLER_51_619 VDD VSS sg13g2_decap_8
XFILLER_63_468 VDD VSS sg13g2_decap_8
XFILLER_90_298 VDD VSS sg13g2_decap_8
XFILLER_32_833 VDD VSS sg13g2_decap_8
XFILLER_17_896 VDD VSS sg13g2_decap_8
XFILLER_31_343 VDD VSS sg13g2_decap_8
X_1713_ _1723_/B _2318_/Q _2304_/Q VDD VSS sg13g2_xnor2_1
XFILLER_99_822 VDD VSS sg13g2_decap_8
X_1644_ _2308_/D VDD _1645_/B VSS _1680_/A _1671_/D sg13g2_o21ai_1
XFILLER_6_84 VDD VSS sg13g2_decap_8
XFILLER_98_332 VDD VSS sg13g2_decap_8
X_1575_ _1575_/Y _1527_/Y _1574_/Y hold484/X _1527_/B VDD VSS sg13g2_a22oi_1
XFILLER_99_866 VDD VSS sg13g2_fill_1
XFILLER_86_505 VDD VSS sg13g2_decap_8
XFILLER_86_549 VDD VSS sg13g2_decap_8
X_2181__178 VDD VSS _2181_/RESET_B sg13g2_tiehi
XFILLER_112_175 VDD VSS sg13g2_decap_8
XFILLER_98_376 VDD VSS sg13g2_decap_8
XFILLER_67_752 VDD VSS sg13g2_fill_1
XFILLER_6_1022 VDD VSS sg13g2_decap_8
XFILLER_39_443 VDD VSS sg13g2_decap_8
XFILLER_55_936 VDD VSS sg13g2_decap_8
XFILLER_27_616 VDD VSS sg13g2_decap_8
XFILLER_66_251 VDD VSS sg13g2_decap_8
XFILLER_82_744 VDD VSS sg13g2_decap_8
XFILLER_81_210 VDD VSS sg13g2_decap_8
X_2127_ _2127_/A _2127_/B _2368_/D VDD VSS sg13g2_nor2_1
XFILLER_54_446 VDD VSS sg13g2_decap_8
XFILLER_26_126 VDD VSS sg13g2_decap_8
X_2058_ _2056_/X _2057_/X _2079_/S _2083_/A VDD VSS sg13g2_mux2_1
XFILLER_70_906 VDD VSS sg13g2_decap_8
XFILLER_82_799 VDD VSS sg13g2_decap_8
XFILLER_81_298 VDD VSS sg13g2_decap_8
XFILLER_63_980 VDD VSS sg13g2_decap_4
XFILLER_35_693 VDD VSS sg13g2_decap_8
XFILLER_23_833 VDD VSS sg13g2_decap_8
XFILLER_25_49 VDD VSS sg13g2_decap_8
XFILLER_22_343 VDD VSS sg13g2_decap_8
XFILLER_50_685 VDD VSS sg13g2_decap_8
XFILLER_109_938 VDD VSS sg13g2_decap_8
XFILLER_108_415 VDD VSS sg13g2_decap_8
XFILLER_89_321 VDD VSS sg13g2_decap_8
Xhold550 _2219_/Q VDD VSS hold550/X sg13g2_dlygate4sd3_1
Xhold561 _2368_/Q VDD VSS hold561/X sg13g2_dlygate4sd3_1
XFILLER_1_203 VDD VSS sg13g2_decap_8
XFILLER_104_654 VDD VSS sg13g2_decap_8
XFILLER_103_175 VDD VSS sg13g2_decap_8
XFILLER_89_398 VDD VSS sg13g2_decap_8
XFILLER_77_516 VDD VSS sg13g2_decap_8
XFILLER_106_63 VDD VSS sg13g2_decap_8
XFILLER_49_207 VDD VSS sg13g2_fill_1
XFILLER_73_700 VDD VSS sg13g2_decap_8
XFILLER_92_519 VDD VSS sg13g2_decap_8
XFILLER_46_925 VDD VSS sg13g2_fill_2
XFILLER_57_262 VDD VSS sg13g2_decap_8
XFILLER_18_616 VDD VSS sg13g2_decap_8
XFILLER_66_56 VDD VSS sg13g2_decap_8
XFILLER_45_402 VDD VSS sg13g2_decap_8
XFILLER_85_582 VDD VSS sg13g2_decap_8
XFILLER_72_221 VDD VSS sg13g2_decap_8
XFILLER_17_126 VDD VSS sg13g2_decap_8
XFILLER_72_243 VDD VSS sg13g2_decap_8
XFILLER_60_405 VDD VSS sg13g2_decap_8
XFILLER_72_287 VDD VSS sg13g2_decap_8
XFILLER_26_693 VDD VSS sg13g2_decap_8
XFILLER_14_833 VDD VSS sg13g2_decap_8
XFILLER_82_77 VDD VSS sg13g2_decap_8
XFILLER_60_449 VDD VSS sg13g2_decap_8
XFILLER_13_343 VDD VSS sg13g2_decap_8
XFILLER_41_685 VDD VSS sg13g2_decap_8
XFILLER_40_140 VDD VSS sg13g2_decap_8
XFILLER_51_1010 VDD VSS sg13g2_decap_8
XFILLER_9_336 VDD VSS sg13g2_decap_8
XFILLER_31_70 VDD VSS sg13g2_decap_8
XFILLER_5_553 VDD VSS sg13g2_decap_8
XFILLER_49_7 VDD VSS sg13g2_decap_8
XFILLER_96_803 VDD VSS sg13g2_fill_1
X_1360_ _1360_/Y _1347_/Y hold417/X _1346_/Y _1385_/A VDD VSS sg13g2_a22oi_1
XFILLER_110_613 VDD VSS sg13g2_decap_8
XFILLER_96_836 VDD VSS sg13g2_decap_8
XFILLER_1_770 VDD VSS sg13g2_decap_8
X_1291_ VDD _2175_/D _1291_/A VSS sg13g2_inv_1
XFILLER_95_357 VDD VSS sg13g2_fill_1
XFILLER_95_335 VDD VSS sg13g2_decap_8
XFILLER_0_280 VDD VSS sg13g2_decap_8
XFILLER_76_571 VDD VSS sg13g2_fill_1
XFILLER_64_711 VDD VSS sg13g2_decap_8
XFILLER_37_903 VDD VSS sg13g2_decap_8
XFILLER_76_582 VDD VSS sg13g2_decap_8
XFILLER_36_413 VDD VSS sg13g2_decap_8
XFILLER_48_295 VDD VSS sg13g2_decap_8
XFILLER_91_563 VDD VSS sg13g2_decap_8
XFILLER_64_788 VDD VSS sg13g2_decap_8
XFILLER_63_243 VDD VSS sg13g2_fill_1
XFILLER_63_276 VDD VSS sg13g2_decap_8
XFILLER_108_1011 VDD VSS sg13g2_decap_8
XFILLER_32_630 VDD VSS sg13g2_decap_8
XFILLER_17_693 VDD VSS sg13g2_decap_8
XFILLER_31_140 VDD VSS sg13g2_decap_8
X_2332__181 VDD VSS _2332_/RESET_B sg13g2_tiehi
XFILLER_20_847 VDD VSS sg13g2_decap_8
XFILLER_75_0 VDD VSS sg13g2_decap_8
X_2367__244 VDD VSS _2367_/RESET_B sg13g2_tiehi
XFILLER_105_407 VDD VSS sg13g2_decap_8
XFILLER_28_1001 VDD VSS sg13g2_decap_8
X_1627_ _1637_/B _2295_/Q _2280_/Q VDD VSS sg13g2_xnor2_1
XFILLER_99_652 VDD VSS sg13g2_decap_8
XFILLER_98_140 VDD VSS sg13g2_decap_8
XFILLER_87_836 VDD VSS sg13g2_decap_8
X_1558_ VSS VDD _1573_/A1 _1211_/Y _1558_/Y _1523_/B sg13g2_a21oi_1
XFILLER_86_335 VDD VSS sg13g2_decap_8
XFILLER_100_112 VDD VSS sg13g2_decap_8
X_1489_ _1236_/C VDD _1497_/A VSS _1235_/A _1234_/B sg13g2_o21ai_1
XFILLER_100_156 VDD VSS sg13g2_fill_1
XFILLER_67_560 VDD VSS sg13g2_decap_8
XFILLER_28_903 VDD VSS sg13g2_decap_8
XFILLER_54_210 VDD VSS sg13g2_decap_4
XFILLER_27_413 VDD VSS sg13g2_decap_8
XFILLER_39_273 VDD VSS sg13g2_decap_8
XFILLER_39_284 VDD VSS sg13g2_fill_2
XFILLER_82_541 VDD VSS sg13g2_decap_8
XFILLER_70_703 VDD VSS sg13g2_decap_8
XFILLER_55_755 VDD VSS sg13g2_decap_8
XFILLER_74_1010 VDD VSS sg13g2_decap_8
XFILLER_36_980 VDD VSS sg13g2_decap_8
XFILLER_42_405 VDD VSS sg13g2_decap_8
XFILLER_23_630 VDD VSS sg13g2_decap_8
XFILLER_52_14 VDD VSS sg13g2_decap_8
XFILLER_35_490 VDD VSS sg13g2_decap_8
XFILLER_22_140 VDD VSS sg13g2_decap_8
XFILLER_52_47 VDD VSS sg13g2_fill_1
XFILLER_11_847 VDD VSS sg13g2_decap_8
XFILLER_52_69 VDD VSS sg13g2_fill_2
XFILLER_10_357 VDD VSS sg13g2_decap_8
XFILLER_109_735 VDD VSS sg13g2_decap_8
XFILLER_108_278 VDD VSS sg13g2_decap_4
XFILLER_105_952 VDD VSS sg13g2_decap_8
XFILLER_89_140 VDD VSS sg13g2_decap_8
Xhold380 _1266_/Y VDD VSS _1267_/A sg13g2_dlygate4sd3_1
XFILLER_104_484 VDD VSS sg13g2_decap_8
XFILLER_104_451 VDD VSS sg13g2_decap_8
Xhold391 _2263_/Q VDD VSS _1485_/A sg13g2_dlygate4sd3_1
XFILLER_2_567 VDD VSS sg13g2_decap_8
XFILLER_77_77 VDD VSS sg13g2_decap_8
XFILLER_93_839 VDD VSS sg13g2_decap_8
XFILLER_92_305 VDD VSS sg13g2_decap_8
XFILLER_65_508 VDD VSS sg13g2_fill_2
XFILLER_19_903 VDD VSS sg13g2_decap_8
XFILLER_93_21 VDD VSS sg13g2_decap_8
XFILLER_46_733 VDD VSS sg13g2_decap_8
XFILLER_18_413 VDD VSS sg13g2_decap_8
XFILLER_45_210 VDD VSS sg13g2_decap_8
XFILLER_73_552 VDD VSS sg13g2_decap_4
XFILLER_85_390 VDD VSS sg13g2_decap_8
XFILLER_34_917 VDD VSS sg13g2_decap_8
XFILLER_45_221 VDD VSS sg13g2_fill_2
XFILLER_73_574 VDD VSS sg13g2_fill_2
XFILLER_93_98 VDD VSS sg13g2_decap_8
XFILLER_27_980 VDD VSS sg13g2_decap_8
XFILLER_61_714 VDD VSS sg13g2_decap_8
XFILLER_33_427 VDD VSS sg13g2_decap_8
XFILLER_60_235 VDD VSS sg13g2_decap_8
XFILLER_14_630 VDD VSS sg13g2_decap_8
XFILLER_26_70 VDD VSS sg13g2_decap_8
XFILLER_26_490 VDD VSS sg13g2_decap_8
XFILLER_13_140 VDD VSS sg13g2_decap_8
XFILLER_42_994 VDD VSS sg13g2_decap_8
XFILLER_9_133 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_6_0 IOVDD IOVSS VDD VSS sg13g2_Filler400
XFILLER_42_91 VDD VSS sg13g2_decap_8
XFILLER_6_840 VDD VSS sg13g2_decap_8
XFILLER_5_350 VDD VSS sg13g2_decap_8
XIO_BOND_iovss_pads\[0\].iovss_pad IOVSS bondpad_70x70
X_1412_ _1412_/Y _1412_/A _1426_/B VDD VSS sg13g2_nand2_1
XFILLER_111_966 VDD VSS sg13g2_decap_8
XFILLER_96_644 VDD VSS sg13g2_decap_8
X_1343_ VDD _2201_/D _1343_/A VSS sg13g2_inv_1
XFILLER_110_410 VDD VSS sg13g2_decap_8
XFILLER_3_63 VDD VSS sg13g2_decap_8
X_1274_ _1274_/Y _1338_/B1 hold322/X _1338_/A2 _2317_/Q VDD VSS sg13g2_a22oi_1
XFILLER_84_828 VDD VSS sg13g2_decap_4
XFILLER_95_154 VDD VSS sg13g2_decap_8
XFILLER_37_700 VDD VSS sg13g2_decap_8
XFILLER_56_519 VDD VSS sg13g2_decap_8
XFILLER_56_508 VDD VSS sg13g2_fill_1
XFILLER_77_891 VDD VSS sg13g2_decap_8
XFILLER_110_487 VDD VSS sg13g2_decap_8
XFILLER_3_1036 VDD VSS sg13g2_decap_8
XFILLER_36_210 VDD VSS sg13g2_decap_8
XFILLER_97_1043 VDD VSS sg13g2_decap_8
XFILLER_92_861 VDD VSS sg13g2_decap_8
XFILLER_25_917 VDD VSS sg13g2_decap_8
XFILLER_37_777 VDD VSS sg13g2_decap_8
XFILLER_64_585 VDD VSS sg13g2_decap_8
XFILLER_18_980 VDD VSS sg13g2_decap_8
XFILLER_24_427 VDD VSS sg13g2_decap_8
XFILLER_36_287 VDD VSS sg13g2_decap_8
XFILLER_51_202 VDD VSS sg13g2_decap_8
XFILLER_91_382 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_16_clk clkbuf_leaf_0_clk/A clkload1/A VDD VSS sg13g2_buf_8
XFILLER_52_758 VDD VSS sg13g2_decap_8
XFILLER_17_490 VDD VSS sg13g2_decap_8
XFILLER_33_994 VDD VSS sg13g2_decap_8
XFILLER_20_644 VDD VSS sg13g2_decap_8
XFILLER_22_28 VDD VSS sg13g2_decap_8
XFILLER_106_727 VDD VSS sg13g2_decap_8
XFILLER_87_644 VDD VSS sg13g2_decap_8
XFILLER_59_324 VDD VSS sg13g2_decap_4
XFILLER_102_977 VDD VSS sg13g2_decap_8
XFILLER_101_465 VDD VSS sg13g2_decap_8
XFILLER_28_700 VDD VSS sg13g2_decap_8
XFILLER_47_14 VDD VSS sg13g2_decap_8
XFILLER_74_338 VDD VSS sg13g2_decap_8
XFILLER_41_1042 VDD VSS sg13g2_decap_8
XFILLER_27_210 VDD VSS sg13g2_decap_8
XFILLER_83_850 VDD VSS sg13g2_decap_8
XFILLER_103_42 VDD VSS sg13g2_decap_8
XFILLER_28_777 VDD VSS sg13g2_decap_8
XFILLER_16_917 VDD VSS sg13g2_decap_8
XFILLER_55_574 VDD VSS sg13g2_decap_8
XFILLER_15_427 VDD VSS sg13g2_decap_8
XFILLER_43_758 VDD VSS sg13g2_decap_8
XFILLER_63_35 VDD VSS sg13g2_decap_8
XFILLER_27_287 VDD VSS sg13g2_decap_8
XFILLER_70_577 VDD VSS sg13g2_decap_8
XFILLER_63_79 VDD VSS sg13g2_fill_1
XFILLER_24_994 VDD VSS sg13g2_decap_8
XFILLER_11_644 VDD VSS sg13g2_decap_8
XFILLER_50_290 VDD VSS sg13g2_decap_8
XFILLER_109_532 VDD VSS sg13g2_decap_8
XFILLER_10_154 VDD VSS sg13g2_decap_8
XFILLER_7_637 VDD VSS sg13g2_decap_8
XFILLER_6_147 VDD VSS sg13g2_decap_8
XFILLER_88_21 VDD VSS sg13g2_decap_8
XFILLER_5_0 VDD VSS sg13g2_decap_8
XFILLER_3_854 VDD VSS sg13g2_decap_8
XFILLER_88_98 VDD VSS sg13g2_decap_8
XFILLER_2_364 VDD VSS sg13g2_decap_8
XFILLER_93_614 VDD VSS sg13g2_decap_8
XFILLER_78_666 VDD VSS sg13g2_decap_4
XFILLER_77_154 VDD VSS sg13g2_decap_8
XFILLER_66_817 VDD VSS sg13g2_decap_8
XFILLER_19_700 VDD VSS sg13g2_decap_8
XFILLER_65_327 VDD VSS sg13g2_fill_2
XFILLER_18_210 VDD VSS sg13g2_decap_8
XFILLER_92_157 VDD VSS sg13g2_decap_8
X_2318__238 VDD VSS _2318_/RESET_B sg13g2_tiehi
XFILLER_34_714 VDD VSS sg13g2_decap_8
XFILLER_19_777 VDD VSS sg13g2_decap_8
XFILLER_37_91 VDD VSS sg13g2_decap_8
XFILLER_73_393 VDD VSS sg13g2_decap_8
XFILLER_61_522 VDD VSS sg13g2_decap_8
XFILLER_18_287 VDD VSS sg13g2_decap_8
XFILLER_33_224 VDD VSS sg13g2_decap_8
XFILLER_57_1060 VDD VSS sg13g2_fill_1
XFILLER_18_1022 VDD VSS sg13g2_decap_8
X_1961_ _1961_/Y _1962_/A _1962_/B VDD VSS sg13g2_nand2_1
XFILLER_30_931 VDD VSS sg13g2_decap_8
XFILLER_42_791 VDD VSS sg13g2_decap_8
XFILLER_15_994 VDD VSS sg13g2_decap_8
XFILLER_105_1036 VDD VSS sg13g2_decap_8
X_1892_ _1892_/B _1892_/A _1892_/X VDD VSS sg13g2_xor2_1
XFILLER_69_600 VDD VSS sg13g2_decap_8
Xclkbuf_leaf_5_clk clkbuf_leaf_5_clk/A clkload7/A VDD VSS sg13g2_buf_8
XFILLER_88_408 VDD VSS sg13g2_decap_8
XFILLER_64_1042 VDD VSS sg13g2_decap_8
XFILLER_25_1015 VDD VSS sg13g2_decap_8
X_2375_ _2375_/RESET_B VSS VDD _2375_/D _2375_/Q clkload8/A sg13g2_dfrbpq_1
XFILLER_38_0 VDD VSS sg13g2_decap_8
XFILLER_68_110 VDD VSS sg13g2_decap_8
XFILLER_111_763 VDD VSS sg13g2_decap_8
X_1326_ _1326_/Y _1342_/B1 hold362/X _1342_/A2 _2326_/Q VDD VSS sg13g2_a22oi_1
XFILLER_96_441 VDD VSS sg13g2_decap_8
XFILLER_57_828 VDD VSS sg13g2_decap_4
XFILLER_56_305 VDD VSS sg13g2_decap_8
XFILLER_112_1029 VDD VSS sg13g2_decap_8
XFILLER_69_699 VDD VSS sg13g2_decap_8
XFILLER_110_273 VDD VSS sg13g2_decap_8
XFILLER_68_176 VDD VSS sg13g2_decap_8
XFILLER_84_669 VDD VSS sg13g2_decap_8
XFILLER_65_850 VDD VSS sg13g2_decap_4
X_1257_ _1257_/Y _1259_/A _1257_/B VDD VSS sg13g2_nand2_1
XFILLER_17_28 VDD VSS sg13g2_decap_8
XFILLER_83_168 VDD VSS sg13g2_decap_4
XFILLER_71_308 VDD VSS sg13g2_decap_8
X_1188_ VDD _2120_/A _1259_/A VSS sg13g2_inv_1
XFILLER_37_574 VDD VSS sg13g2_decap_8
XFILLER_25_714 VDD VSS sg13g2_decap_8
XFILLER_52_533 VDD VSS sg13g2_decap_8
XFILLER_24_224 VDD VSS sg13g2_decap_8
XFILLER_52_555 VDD VSS sg13g2_decap_8
XFILLER_21_931 VDD VSS sg13g2_decap_8
XFILLER_40_739 VDD VSS sg13g2_decap_8
XFILLER_33_791 VDD VSS sg13g2_decap_8
XFILLER_33_49 VDD VSS sg13g2_decap_8
XFILLER_32_1008 VDD VSS sg13g2_decap_8
XFILLER_20_441 VDD VSS sg13g2_decap_8
XFILLER_79_419 VDD VSS sg13g2_decap_8
XFILLER_99_290 VDD VSS sg13g2_decap_8
XFILLER_87_430 VDD VSS sg13g2_decap_8
XFILLER_59_110 VDD VSS sg13g2_decap_8
XFILLER_88_986 VDD VSS sg13g2_decap_8
XFILLER_102_752 VDD VSS sg13g2_decap_4
XFILLER_48_828 VDD VSS sg13g2_decap_8
XFILLER_0_868 VDD VSS sg13g2_decap_8
XFILLER_58_79 VDD VSS sg13g2_decap_8
XFILLER_101_262 VDD VSS sg13g2_decap_8
XFILLER_47_338 VDD VSS sg13g2_decap_8
XFILLER_75_658 VDD VSS sg13g2_decap_8
XFILLER_56_850 VDD VSS sg13g2_decap_8
XFILLER_74_56 VDD VSS sg13g2_decap_8
XFILLER_28_574 VDD VSS sg13g2_decap_8
XFILLER_16_714 VDD VSS sg13g2_decap_8
X_2303__99 VDD VSS _2303__99/L_HI sg13g2_tiehi
XFILLER_83_691 VDD VSS sg13g2_decap_8
XFILLER_15_224 VDD VSS sg13g2_decap_8
XFILLER_70_341 VDD VSS sg13g2_fill_1
XFILLER_31_728 VDD VSS sg13g2_decap_8
XFILLER_24_791 VDD VSS sg13g2_decap_8
XFILLER_12_931 VDD VSS sg13g2_decap_8
XFILLER_90_77 VDD VSS sg13g2_decap_8
XFILLER_11_441 VDD VSS sg13g2_decap_8
XFILLER_30_238 VDD VSS sg13g2_decap_8
XFILLER_8_924 VDD VSS sg13g2_decap_8
XFILLER_109_340 VDD VSS sg13g2_decap_8
XFILLER_7_434 VDD VSS sg13g2_decap_8
XFILLER_99_42 VDD VSS sg13g2_decap_8
XFILLER_79_920 VDD VSS sg13g2_decap_8
XFILLER_48_1037 VDD VSS sg13g2_decap_8
XFILLER_3_651 VDD VSS sg13g2_decap_8
XFILLER_97_249 VDD VSS sg13g2_decap_8
XFILLER_2_161 VDD VSS sg13g2_decap_8
XFILLER_31_7 VDD VSS sg13g2_decap_8
XFILLER_79_975 VDD VSS sg13g2_decap_8
XFILLER_94_934 VDD VSS sg13g2_decap_8
X_2160_ _2162_/A _2160_/B _2348_/D VDD VSS sg13g2_nor2_1
XFILLER_78_485 VDD VSS sg13g2_decap_4
XFILLER_38_327 VDD VSS sg13g2_decap_8
X_2091_ _2162_/A _2156_/A _2344_/D VDD VSS sg13g2_nor2_1
XFILLER_80_105 VDD VSS sg13g2_decap_8
XFILLER_0_42 VDD VSS sg13g2_decap_8
XFILLER_19_574 VDD VSS sg13g2_decap_8
XFILLER_47_894 VDD VSS sg13g2_decap_8
XFILLER_34_511 VDD VSS sg13g2_decap_8
XFILLER_46_393 VDD VSS sg13g2_decap_8
XFILLER_62_864 VDD VSS sg13g2_decap_8
XFILLER_34_588 VDD VSS sg13g2_decap_8
XFILLER_22_728 VDD VSS sg13g2_decap_8
XFILLER_15_791 VDD VSS sg13g2_decap_8
X_1944_ _1938_/B _1938_/A _1932_/Y _1946_/B VDD VSS sg13g2_a21o_1
XFILLER_21_238 VDD VSS sg13g2_decap_8
XFILLER_9_84 VDD VSS sg13g2_decap_8
X_1875_ _1876_/B _1884_/A _1884_/B VDD VSS sg13g2_nand2b_1
XFILLER_89_706 VDD VSS sg13g2_decap_8
XFILLER_97_750 VDD VSS sg13g2_decap_8
XFILLER_111_560 VDD VSS sg13g2_decap_8
XFILLER_57_625 VDD VSS sg13g2_decap_8
X_2358_ _2358_/RESET_B VSS VDD _2358_/D _2358_/Q clkload2/A sg13g2_dfrbpq_1
X_1309_ VDD _2184_/D _1309_/A VSS sg13g2_inv_1
XFILLER_28_49 VDD VSS sg13g2_decap_8
XFILLER_56_124 VDD VSS sg13g2_decap_8
X_2289_ _2289_/RESET_B VSS VDD _2289_/D _2289_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_84_466 VDD VSS sg13g2_decap_8
XFILLER_44_308 VDD VSS sg13g2_decap_8
XFILLER_71_138 VDD VSS sg13g2_fill_1
XFILLER_53_831 VDD VSS sg13g2_decap_8
XFILLER_25_511 VDD VSS sg13g2_decap_8
XFILLER_37_371 VDD VSS sg13g2_decap_8
XFILLER_52_341 VDD VSS sg13g2_decap_4
XFILLER_52_352 VDD VSS sg13g2_decap_8
X_2191__158 VDD VSS _2191_/RESET_B sg13g2_tiehi
XFILLER_100_21 VDD VSS sg13g2_decap_8
XFILLER_25_588 VDD VSS sg13g2_decap_8
XFILLER_52_396 VDD VSS sg13g2_decap_8
XFILLER_13_728 VDD VSS sg13g2_decap_8
XFILLER_12_238 VDD VSS sg13g2_decap_8
XFILLER_100_98 VDD VSS sg13g2_decap_8
XFILLER_60_14 VDD VSS sg13g2_decap_8
XFILLER_60_25 VDD VSS sg13g2_fill_2
XFILLER_107_800 VDD VSS sg13g2_decap_8
XFILLER_5_938 VDD VSS sg13g2_decap_8
XFILLER_109_63 VDD VSS sg13g2_decap_8
XFILLER_4_448 VDD VSS sg13g2_decap_8
XFILLER_107_877 VDD VSS sg13g2_decap_8
XFILLER_106_365 VDD VSS sg13g2_decap_8
X_2221__98 VDD VSS _2221__98/L_HI sg13g2_tiehi
XFILLER_88_761 VDD VSS sg13g2_fill_2
XFILLER_88_750 VDD VSS sg13g2_decap_8
XFILLER_48_603 VDD VSS sg13g2_decap_8
XFILLER_0_665 VDD VSS sg13g2_decap_8
XFILLER_75_411 VDD VSS sg13g2_decap_8
XFILLER_85_77 VDD VSS sg13g2_decap_8
XFILLER_47_146 VDD VSS sg13g2_fill_2
XFILLER_91_926 VDD VSS sg13g2_decap_8
XFILLER_78_1008 VDD VSS sg13g2_fill_2
XFILLER_63_628 VDD VSS sg13g2_decap_8
XFILLER_29_861 VDD VSS sg13g2_decap_8
XFILLER_62_105 VDD VSS sg13g2_decap_8
XFILLER_35_308 VDD VSS sg13g2_decap_8
XFILLER_44_842 VDD VSS sg13g2_decap_4
XFILLER_16_511 VDD VSS sg13g2_decap_8
XFILLER_62_127 VDD VSS sg13g2_decap_8
XFILLER_28_371 VDD VSS sg13g2_decap_8
XFILLER_71_661 VDD VSS sg13g2_decap_8
XFILLER_90_469 VDD VSS sg13g2_decap_8
XFILLER_71_694 VDD VSS sg13g2_fill_1
XFILLER_44_886 VDD VSS sg13g2_decap_8
XFILLER_16_588 VDD VSS sg13g2_decap_8
XFILLER_31_525 VDD VSS sg13g2_decap_8
XFILLER_43_385 VDD VSS sg13g2_decap_8
XFILLER_70_182 VDD VSS sg13g2_decap_4
XFILLER_34_70 VDD VSS sg13g2_decap_8
XFILLER_8_721 VDD VSS sg13g2_decap_8
XFILLER_15_1036 VDD VSS sg13g2_decap_8
XFILLER_79_7 VDD VSS sg13g2_decap_8
XFILLER_7_231 VDD VSS sg13g2_decap_8
X_1660_ _1660_/Y _1646_/Y _1659_/X hold453/X _1671_/B VDD VSS sg13g2_a22oi_1
XFILLER_8_798 VDD VSS sg13g2_decap_8
X_1591_ _1592_/A _1592_/B _1593_/B VDD VSS sg13g2_nor2_1
XFILLER_98_525 VDD VSS sg13g2_decap_8
XFILLER_79_750 VDD VSS sg13g2_decap_8
XFILLER_112_357 VDD VSS sg13g2_decap_8
XFILLER_61_1012 VDD VSS sg13g2_decap_8
XFILLER_94_720 VDD VSS sg13g2_decap_8
X_2212_ _2212_/RESET_B VSS VDD _2212_/D _2212_/Q _2245_/CLK sg13g2_dfrbpq_1
X_2143_ _2143_/A _2143_/B _2372_/D VDD VSS sg13g2_nor2_1
XFILLER_67_978 VDD VSS sg13g2_decap_8
XFILLER_22_1029 VDD VSS sg13g2_decap_8
XFILLER_39_647 VDD VSS sg13g2_decap_8
XFILLER_94_786 VDD VSS sg13g2_fill_2
XFILLER_54_628 VDD VSS sg13g2_decap_4
XFILLER_26_308 VDD VSS sg13g2_decap_8
XFILLER_38_168 VDD VSS sg13g2_decap_8
X_2074_ _2074_/Y _2074_/A _2074_/B VDD VSS sg13g2_nand2_1
XFILLER_93_296 VDD VSS sg13g2_decap_8
XFILLER_81_447 VDD VSS sg13g2_decap_8
XFILLER_47_691 VDD VSS sg13g2_decap_8
XFILLER_19_371 VDD VSS sg13g2_decap_8
Xin_data_pads\[7\].in_data_pad IOVDD IOVSS _1388_/A in_data_PADs[7] VDD VSS sg13g2_IOPadIn
XFILLER_35_875 VDD VSS sg13g2_decap_8
XFILLER_50_812 VDD VSS sg13g2_decap_8
XFILLER_61_171 VDD VSS sg13g2_decap_8
XFILLER_22_525 VDD VSS sg13g2_decap_8
XFILLER_34_385 VDD VSS sg13g2_decap_8
X_1927_ _1927_/A _1940_/A _1928_/B VDD VSS sg13g2_nor2_1
XFILLER_108_619 VDD VSS sg13g2_decap_8
X_1858_ _2203_/Q _2244_/Q _2048_/A VDD VSS sg13g2_xor2_1
XFILLER_30_28 VDD VSS sg13g2_decap_8
Xfanout3 _2043_/S _2089_/S VDD VSS sg13g2_buf_1
X_1789_ VDD VSS _1817_/B _1778_/Y _1900_/A _1777_/Y _1812_/A _1779_/Y sg13g2_a221oi_1
XFILLER_103_313 VDD VSS sg13g2_decap_8
XFILLER_89_558 VDD VSS sg13g2_decap_8
XFILLER_77_709 VDD VSS sg13g2_decap_8
XFILLER_58_901 VDD VSS sg13g2_decap_8
XFILLER_76_219 VDD VSS sg13g2_decap_8
XFILLER_69_260 VDD VSS sg13g2_decap_8
XFILLER_57_411 VDD VSS sg13g2_decap_8
XFILLER_97_591 VDD VSS sg13g2_fill_2
XFILLER_85_742 VDD VSS sg13g2_decap_8
XFILLER_73_915 VDD VSS sg13g2_decap_4
XFILLER_84_241 VDD VSS sg13g2_decap_8
XFILLER_17_308 VDD VSS sg13g2_decap_8
XFILLER_55_14 VDD VSS sg13g2_decap_8
XFILLER_29_168 VDD VSS sg13g2_decap_8
XFILLER_84_285 VDD VSS sg13g2_decap_8
XFILLER_72_414 VDD VSS sg13g2_decap_8
XFILLER_72_425 VDD VSS sg13g2_fill_1
XFILLER_44_127 VDD VSS sg13g2_decap_8
XFILLER_72_469 VDD VSS sg13g2_decap_8
XFILLER_38_1003 VDD VSS sg13g2_decap_8
XFILLER_26_875 VDD VSS sg13g2_decap_8
XFILLER_81_981 VDD VSS sg13g2_fill_2
XFILLER_111_42 VDD VSS sg13g2_decap_8
XFILLER_53_683 VDD VSS sg13g2_decap_8
XFILLER_13_525 VDD VSS sg13g2_decap_8
XFILLER_25_385 VDD VSS sg13g2_decap_8
XFILLER_40_300 VDD VSS sg13g2_decap_8
XFILLER_52_171 VDD VSS sg13g2_fill_1
XFILLER_71_35 VDD VSS sg13g2_decap_8
XFILLER_41_867 VDD VSS sg13g2_decap_8
X_2314__263 VDD VSS _2314_/RESET_B sg13g2_tiehi
XFILLER_9_518 VDD VSS sg13g2_decap_8
XFILLER_40_377 VDD VSS sg13g2_decap_8
XFILLER_5_735 VDD VSS sg13g2_decap_8
XFILLER_84_1001 VDD VSS sg13g2_decap_8
XFILLER_84_1023 VDD VSS sg13g2_decap_8
XFILLER_107_674 VDD VSS sg13g2_decap_8
XFILLER_106_140 VDD VSS sg13g2_decap_8
XFILLER_105_0 VDD VSS sg13g2_decap_8
XFILLER_4_245 VDD VSS sg13g2_decap_8
XFILLER_96_21 VDD VSS sg13g2_decap_8
XFILLER_1_952 VDD VSS sg13g2_decap_8
XFILLER_76_720 VDD VSS sg13g2_decap_8
XFILLER_0_462 VDD VSS sg13g2_decap_8
XFILLER_96_98 VDD VSS sg13g2_decap_8
XFILLER_49_945 VDD VSS sg13g2_fill_2
XFILLER_29_70 VDD VSS sg13g2_decap_8
XFILLER_48_444 VDD VSS sg13g2_decap_8
XFILLER_64_915 VDD VSS sg13g2_fill_1
XFILLER_91_745 VDD VSS sg13g2_decap_8
XFILLER_76_797 VDD VSS sg13g2_decap_8
XFILLER_75_285 VDD VSS sg13g2_decap_8
XFILLER_63_447 VDD VSS sg13g2_decap_8
XFILLER_35_105 VDD VSS sg13g2_decap_8
XFILLER_17_875 VDD VSS sg13g2_decap_8
XFILLER_90_277 VDD VSS sg13g2_decap_8
XFILLER_90_288 VDD VSS sg13g2_fill_1
XFILLER_44_683 VDD VSS sg13g2_decap_8
XFILLER_32_812 VDD VSS sg13g2_decap_8
XFILLER_16_385 VDD VSS sg13g2_decap_8
XFILLER_45_91 VDD VSS sg13g2_decap_4
XFILLER_91_1049 VDD VSS sg13g2_decap_8
XFILLER_31_322 VDD VSS sg13g2_decap_8
XFILLER_43_182 VDD VSS sg13g2_decap_8
XFILLER_32_889 VDD VSS sg13g2_decap_8
XFILLER_31_399 VDD VSS sg13g2_decap_8
X_1712_ _1725_/A _1712_/B _1712_/Y VDD VSS sg13g2_nor2_1
XFILLER_61_90 VDD VSS sg13g2_decap_8
X_1643_ _1671_/B _1671_/C _2308_/D VDD VSS sg13g2_nor2_1
XFILLER_8_595 VDD VSS sg13g2_decap_8
XFILLER_99_801 VDD VSS sg13g2_decap_8
XFILLER_6_63 VDD VSS sg13g2_decap_8
X_1574_ _1573_/Y VDD _1574_/Y VSS _2288_/Q _1571_/Y sg13g2_o21ai_1
XIO_FILL_IO_EAST_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_99_889 VDD VSS sg13g2_fill_1
XFILLER_101_828 VDD VSS sg13g2_decap_8
XFILLER_86_517 VDD VSS sg13g2_decap_8
XFILLER_112_154 VDD VSS sg13g2_decap_8
XFILLER_58_208 VDD VSS sg13g2_decap_8
XFILLER_6_1001 VDD VSS sg13g2_decap_8
XFILLER_100_349 VDD VSS sg13g2_decap_8
XFILLER_20_0 VDD VSS sg13g2_decap_8
XFILLER_39_422 VDD VSS sg13g2_decap_8
XFILLER_66_230 VDD VSS sg13g2_decap_4
XFILLER_94_594 VDD VSS sg13g2_decap_8
XFILLER_82_723 VDD VSS sg13g2_decap_8
X_2126_ _1688_/B VDD _2127_/B VSS _1259_/A hold561/X sg13g2_o21ai_1
XFILLER_55_959 VDD VSS sg13g2_decap_8
XFILLER_54_425 VDD VSS sg13g2_decap_8
XFILLER_26_105 VDD VSS sg13g2_decap_8
XFILLER_39_499 VDD VSS sg13g2_decap_8
XFILLER_82_778 VDD VSS sg13g2_decap_8
X_2057_ _1953_/A _1892_/X _2069_/S _2057_/X VDD VSS sg13g2_mux2_1
XFILLER_42_609 VDD VSS sg13g2_decap_8
XFILLER_81_277 VDD VSS sg13g2_decap_8
XFILLER_35_672 VDD VSS sg13g2_decap_8
XFILLER_23_812 VDD VSS sg13g2_decap_8
XFILLER_25_28 VDD VSS sg13g2_decap_8
XFILLER_41_119 VDD VSS sg13g2_decap_8
XFILLER_62_491 VDD VSS sg13g2_decap_8
XFILLER_22_322 VDD VSS sg13g2_decap_8
XFILLER_34_182 VDD VSS sg13g2_decap_8
XFILLER_50_664 VDD VSS sg13g2_decap_8
XFILLER_23_889 VDD VSS sg13g2_decap_8
XFILLER_10_539 VDD VSS sg13g2_decap_8
XFILLER_22_399 VDD VSS sg13g2_decap_8
XFILLER_109_917 VDD VSS sg13g2_decap_8
XFILLER_41_49 VDD VSS sg13g2_decap_8
XIO_BOND_iovdd_pads\[0\].iovdd_pad IOVDD bondpad_70x70
Xhold540 _1717_/Y VDD VSS _1718_/B sg13g2_dlygate4sd3_1
XFILLER_89_300 VDD VSS sg13g2_decap_8
XFILLER_9_7 VDD VSS sg13g2_decap_8
XFILLER_2_749 VDD VSS sg13g2_decap_8
Xhold562 _2283_/Q VDD VSS hold562/X sg13g2_dlygate4sd3_1
Xhold551 _2293_/Q VDD VSS hold551/X sg13g2_dlygate4sd3_1
XFILLER_104_633 VDD VSS sg13g2_decap_8
XFILLER_1_259 VDD VSS sg13g2_decap_8
XFILLER_89_377 VDD VSS sg13g2_decap_8
XFILLER_106_42 VDD VSS sg13g2_decap_8
XFILLER_103_154 VDD VSS sg13g2_decap_8
XFILLER_44_1040 VDD VSS sg13g2_decap_8
XFILLER_49_219 VDD VSS sg13g2_fill_2
XFILLER_58_742 VDD VSS sg13g2_decap_8
XFILLER_58_753 VDD VSS sg13g2_fill_1
XFILLER_66_35 VDD VSS sg13g2_decap_8
XFILLER_100_861 VDD VSS sg13g2_decap_8
XFILLER_85_561 VDD VSS sg13g2_decap_8
XFILLER_46_904 VDD VSS sg13g2_decap_8
XFILLER_17_105 VDD VSS sg13g2_decap_8
XFILLER_45_414 VDD VSS sg13g2_decap_8
XFILLER_33_609 VDD VSS sg13g2_decap_8
XFILLER_45_469 VDD VSS sg13g2_decap_8
XFILLER_73_789 VDD VSS sg13g2_decap_8
XFILLER_82_56 VDD VSS sg13g2_decap_8
XFILLER_26_672 VDD VSS sg13g2_decap_8
XFILLER_14_812 VDD VSS sg13g2_decap_8
XFILLER_32_119 VDD VSS sg13g2_decap_8
XFILLER_53_491 VDD VSS sg13g2_decap_8
XFILLER_13_322 VDD VSS sg13g2_decap_8
XFILLER_25_182 VDD VSS sg13g2_decap_8
XFILLER_41_664 VDD VSS sg13g2_decap_8
XFILLER_9_315 VDD VSS sg13g2_decap_8
XFILLER_14_889 VDD VSS sg13g2_decap_8
XFILLER_13_399 VDD VSS sg13g2_decap_8
XFILLER_40_196 VDD VSS sg13g2_decap_8
XFILLER_5_532 VDD VSS sg13g2_decap_8
XIO_BOND_out_data_pads\[0\].out_data_pad out_data_PADs[0] bondpad_70x70
XFILLER_108_983 VDD VSS sg13g2_decap_8
XFILLER_99_119 VDD VSS sg13g2_decap_8
XFILLER_96_815 VDD VSS sg13g2_decap_8
XFILLER_95_314 VDD VSS sg13g2_decap_8
X_1290_ _1290_/Y _1322_/B1 hold360/X _1322_/A2 _2339_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_669 VDD VSS sg13g2_decap_8
XFILLER_48_230 VDD VSS sg13g2_decap_8
XFILLER_37_959 VDD VSS sg13g2_decap_8
XFILLER_49_797 VDD VSS sg13g2_decap_8
X_2351__97 VDD VSS _2351__97/L_HI sg13g2_tiehi
XFILLER_48_274 VDD VSS sg13g2_decap_8
XFILLER_91_542 VDD VSS sg13g2_decap_8
XFILLER_64_767 VDD VSS sg13g2_decap_8
XFILLER_24_609 VDD VSS sg13g2_decap_8
XFILLER_63_255 VDD VSS sg13g2_decap_8
XFILLER_36_469 VDD VSS sg13g2_decap_8
XFILLER_52_929 VDD VSS sg13g2_decap_8
XFILLER_51_406 VDD VSS sg13g2_fill_2
XFILLER_17_672 VDD VSS sg13g2_decap_8
XFILLER_23_119 VDD VSS sg13g2_decap_8
XFILLER_16_182 VDD VSS sg13g2_decap_8
XFILLER_32_686 VDD VSS sg13g2_decap_8
XFILLER_20_826 VDD VSS sg13g2_decap_8
XFILLER_31_196 VDD VSS sg13g2_decap_8
XFILLER_9_882 VDD VSS sg13g2_decap_8
XFILLER_68_0 VDD VSS sg13g2_decap_8
XFILLER_106_909 VDD VSS sg13g2_decap_8
XFILLER_8_392 VDD VSS sg13g2_decap_8
X_1626_ _1639_/A _1626_/B _1626_/Y VDD VSS sg13g2_nor2_1
X_1557_ VDD _1557_/Y _1557_/A VSS sg13g2_inv_1
XFILLER_87_815 VDD VSS sg13g2_decap_8
XFILLER_86_314 VDD VSS sg13g2_decap_8
XFILLER_28_1057 VDD VSS sg13g2_decap_4
XFILLER_101_636 VDD VSS sg13g2_decap_8
XFILLER_59_539 VDD VSS sg13g2_decap_8
X_1488_ VSS VDD _1252_/Y hold341/X _1488_/Y _2101_/A sg13g2_a21oi_1
XFILLER_39_252 VDD VSS sg13g2_decap_8
XFILLER_82_520 VDD VSS sg13g2_decap_8
XFILLER_28_959 VDD VSS sg13g2_decap_8
XFILLER_55_734 VDD VSS sg13g2_decap_8
XFILLER_94_391 VDD VSS sg13g2_decap_8
X_2109_ _1510_/A _2195_/Q _2187_/Q _2179_/Q _2171_/Q _1510_/B _2109_/X VDD VSS sg13g2_mux4_1
XFILLER_55_778 VDD VSS sg13g2_fill_1
XFILLER_15_609 VDD VSS sg13g2_decap_8
XFILLER_36_49 VDD VSS sg13g2_decap_8
XFILLER_27_469 VDD VSS sg13g2_decap_8
XFILLER_82_597 VDD VSS sg13g2_fill_2
XFILLER_14_119 VDD VSS sg13g2_decap_8
XFILLER_70_759 VDD VSS sg13g2_decap_8
X_2270__214 VDD VSS _2270_/RESET_B sg13g2_tiehi
XFILLER_54_299 VDD VSS sg13g2_decap_8
XFILLER_23_686 VDD VSS sg13g2_decap_8
XFILLER_11_826 VDD VSS sg13g2_decap_8
XFILLER_50_472 VDD VSS sg13g2_decap_8
XFILLER_109_714 VDD VSS sg13g2_decap_8
XFILLER_10_336 VDD VSS sg13g2_decap_8
XFILLER_7_819 VDD VSS sg13g2_decap_8
XFILLER_22_196 VDD VSS sg13g2_decap_8
XFILLER_6_329 VDD VSS sg13g2_decap_8
XFILLER_108_257 VDD VSS sg13g2_decap_8
XFILLER_11_1050 VDD VSS sg13g2_decap_8
XFILLER_105_931 VDD VSS sg13g2_decap_8
Xhold381 _2194_/Q VDD VSS hold381/X sg13g2_dlygate4sd3_1
XFILLER_104_430 VDD VSS sg13g2_decap_8
Xhold370 _2252_/Q VDD VSS _1201_/A sg13g2_dlygate4sd3_1
XFILLER_2_546 VDD VSS sg13g2_decap_8
XFILLER_81_1015 VDD VSS sg13g2_decap_8
Xhold392 _1485_/Y VDD VSS hold392/X sg13g2_dlygate4sd3_1
XFILLER_81_1059 VDD VSS sg13g2_fill_2
XFILLER_81_1048 VDD VSS sg13g2_decap_8
XFILLER_77_336 VDD VSS sg13g2_decap_8
XFILLER_77_56 VDD VSS sg13g2_decap_8
XFILLER_93_818 VDD VSS sg13g2_decap_8
XFILLER_19_959 VDD VSS sg13g2_decap_8
XFILLER_73_531 VDD VSS sg13g2_decap_8
XFILLER_18_469 VDD VSS sg13g2_decap_8
XFILLER_73_586 VDD VSS sg13g2_decap_8
XFILLER_93_77 VDD VSS sg13g2_decap_8
XFILLER_61_737 VDD VSS sg13g2_fill_1
XFILLER_46_789 VDD VSS sg13g2_decap_8
XFILLER_33_406 VDD VSS sg13g2_decap_8
XFILLER_60_214 VDD VSS sg13g2_decap_8
XFILLER_42_973 VDD VSS sg13g2_decap_8
XFILLER_9_112 VDD VSS sg13g2_decap_8
XFILLER_14_686 VDD VSS sg13g2_decap_8
XFILLER_13_196 VDD VSS sg13g2_decap_8
XFILLER_42_70 VDD VSS sg13g2_decap_8
XFILLER_9_189 VDD VSS sg13g2_decap_8
XFILLER_61_7 VDD VSS sg13g2_decap_8
XFILLER_108_780 VDD VSS sg13g2_decap_8
XFILLER_6_896 VDD VSS sg13g2_decap_8
X_1411_ VSS VDD _2265_/Q _1410_/B _1426_/B _1429_/A sg13g2_a21oi_1
XFILLER_69_837 VDD VSS sg13g2_fill_2
XFILLER_69_804 VDD VSS sg13g2_fill_1
XFILLER_111_945 VDD VSS sg13g2_decap_8
XFILLER_96_623 VDD VSS sg13g2_decap_8
X_1342_ _1342_/Y _1342_/B1 hold316/X _1342_/A2 _2334_/Q VDD VSS sg13g2_a22oi_1
XFILLER_68_347 VDD VSS sg13g2_decap_8
XFILLER_3_42 VDD VSS sg13g2_decap_8
X_1273_ VDD _2166_/D _1273_/A VSS sg13g2_inv_1
XFILLER_77_870 VDD VSS sg13g2_decap_8
XFILLER_110_466 VDD VSS sg13g2_decap_8
XFILLER_83_306 VDD VSS sg13g2_fill_2
XFILLER_95_133 VDD VSS sg13g2_decap_8
XFILLER_68_369 VDD VSS sg13g2_fill_2
XFILLER_83_339 VDD VSS sg13g2_decap_8
XFILLER_49_572 VDD VSS sg13g2_decap_8
XFILLER_3_1015 VDD VSS sg13g2_decap_8
XFILLER_92_840 VDD VSS sg13g2_decap_8
XFILLER_76_380 VDD VSS sg13g2_decap_8
XFILLER_37_756 VDD VSS sg13g2_decap_8
XFILLER_64_564 VDD VSS sg13g2_decap_8
XFILLER_52_726 VDD VSS sg13g2_decap_4
XFILLER_24_406 VDD VSS sg13g2_decap_8
XFILLER_36_266 VDD VSS sg13g2_decap_8
XFILLER_33_973 VDD VSS sg13g2_decap_8
XFILLER_51_258 VDD VSS sg13g2_decap_8
XFILLER_60_792 VDD VSS sg13g2_decap_8
XFILLER_20_623 VDD VSS sg13g2_decap_8
XFILLER_32_483 VDD VSS sg13g2_decap_8
XFILLER_34_1050 VDD VSS sg13g2_decap_8
XFILLER_106_706 VDD VSS sg13g2_decap_8
XFILLER_105_249 VDD VSS sg13g2_decap_8
Xiovss_pads\[0\].iovss_pad IOVDD IOVSS VDD VSS sg13g2_IOPadIOVss
X_1609_ _1608_/Y VDD _1610_/B VSS _1638_/S hold523/X sg13g2_o21ai_1
XFILLER_102_956 VDD VSS sg13g2_decap_8
XFILLER_87_623 VDD VSS sg13g2_decap_8
XFILLER_101_400 VDD VSS sg13g2_decap_8
XFILLER_99_483 VDD VSS sg13g2_decap_8
XFILLER_87_689 VDD VSS sg13g2_decap_8
XFILLER_101_444 VDD VSS sg13g2_decap_8
XFILLER_41_1021 VDD VSS sg13g2_decap_8
XFILLER_59_369 VDD VSS sg13g2_decap_8
XFILLER_47_509 VDD VSS sg13g2_decap_8
XFILLER_101_499 VDD VSS sg13g2_decap_8
XFILLER_86_199 VDD VSS sg13g2_decap_4
XFILLER_74_328 VDD VSS sg13g2_decap_8
XFILLER_103_21 VDD VSS sg13g2_decap_8
XFILLER_55_553 VDD VSS sg13g2_decap_8
XFILLER_28_756 VDD VSS sg13g2_decap_8
XFILLER_82_361 VDD VSS sg13g2_decap_8
XFILLER_70_512 VDD VSS sg13g2_decap_4
XFILLER_15_406 VDD VSS sg13g2_decap_8
XFILLER_63_14 VDD VSS sg13g2_decap_8
XFILLER_27_266 VDD VSS sg13g2_decap_8
XFILLER_82_394 VDD VSS sg13g2_decap_8
XFILLER_103_98 VDD VSS sg13g2_decap_8
XFILLER_55_597 VDD VSS sg13g2_fill_1
XFILLER_43_737 VDD VSS sg13g2_decap_8
XFILLER_70_556 VDD VSS sg13g2_decap_8
XFILLER_24_973 VDD VSS sg13g2_decap_8
XFILLER_11_623 VDD VSS sg13g2_decap_8
XFILLER_23_483 VDD VSS sg13g2_decap_8
XFILLER_10_133 VDD VSS sg13g2_decap_8
XFILLER_7_616 VDD VSS sg13g2_decap_8
XFILLER_109_511 VDD VSS sg13g2_decap_8
XFILLER_6_126 VDD VSS sg13g2_decap_8
XFILLER_109_588 VDD VSS sg13g2_decap_8
XFILLER_12_84 VDD VSS sg13g2_decap_8
XFILLER_3_833 VDD VSS sg13g2_decap_8
XFILLER_88_77 VDD VSS sg13g2_decap_8
XFILLER_2_343 VDD VSS sg13g2_decap_8
XFILLER_77_133 VDD VSS sg13g2_decap_8
XFILLER_38_509 VDD VSS sg13g2_decap_8
XFILLER_19_756 VDD VSS sg13g2_decap_8
XFILLER_46_531 VDD VSS sg13g2_fill_2
XFILLER_74_873 VDD VSS sg13g2_fill_2
XFILLER_74_884 VDD VSS sg13g2_decap_8
XFILLER_18_266 VDD VSS sg13g2_decap_8
XFILLER_37_70 VDD VSS sg13g2_decap_8
XFILLER_33_203 VDD VSS sg13g2_decap_8
XFILLER_73_372 VDD VSS sg13g2_decap_8
XFILLER_15_973 VDD VSS sg13g2_decap_8
XFILLER_18_1001 VDD VSS sg13g2_decap_8
X_1960_ _1960_/B _1960_/A _1962_/B VDD VSS sg13g2_xor2_1
XFILLER_42_770 VDD VSS sg13g2_decap_8
XFILLER_30_910 VDD VSS sg13g2_decap_8
XFILLER_14_483 VDD VSS sg13g2_decap_8
XFILLER_105_1015 VDD VSS sg13g2_decap_8
X_1891_ _1891_/B _1891_/A _1960_/A VDD VSS sg13g2_xor2_1
XFILLER_30_987 VDD VSS sg13g2_decap_8
XFILLER_6_693 VDD VSS sg13g2_decap_8
XFILLER_64_1021 VDD VSS sg13g2_decap_8
XFILLER_102_219 VDD VSS sg13g2_decap_4
XFILLER_96_420 VDD VSS sg13g2_decap_8
X_2374_ _2374_/RESET_B VSS VDD _2374_/D _2374_/Q clkload1/A sg13g2_dfrbpq_1
XFILLER_111_742 VDD VSS sg13g2_decap_8
X_1325_ VDD _2192_/D _1325_/A VSS sg13g2_inv_1
XFILLER_69_678 VDD VSS sg13g2_decap_8
XFILLER_69_656 VDD VSS sg13g2_decap_8
XFILLER_57_807 VDD VSS sg13g2_decap_8
XFILLER_112_1008 VDD VSS sg13g2_decap_8
XFILLER_97_998 VDD VSS sg13g2_decap_8
XFILLER_110_252 VDD VSS sg13g2_decap_8
XFILLER_96_486 VDD VSS sg13g2_decap_8
XFILLER_84_648 VDD VSS sg13g2_decap_8
XFILLER_83_147 VDD VSS sg13g2_decap_8
X_1256_ _1259_/C _1507_/A _2273_/Q _1257_/B VDD VSS sg13g2_nand3_1
XFILLER_49_391 VDD VSS sg13g2_decap_8
XFILLER_37_553 VDD VSS sg13g2_decap_8
XFILLER_80_832 VDD VSS sg13g2_decap_8
XFILLER_65_895 VDD VSS sg13g2_decap_8
XFILLER_52_512 VDD VSS sg13g2_decap_8
XFILLER_24_203 VDD VSS sg13g2_decap_8
XFILLER_80_887 VDD VSS sg13g2_decap_8
XFILLER_40_718 VDD VSS sg13g2_decap_8
XFILLER_33_770 VDD VSS sg13g2_decap_8
XFILLER_21_910 VDD VSS sg13g2_decap_8
XFILLER_33_28 VDD VSS sg13g2_decap_8
XFILLER_71_1047 VDD VSS sg13g2_decap_8
XFILLER_20_420 VDD VSS sg13g2_decap_8
XFILLER_32_280 VDD VSS sg13g2_decap_8
XFILLER_21_987 VDD VSS sg13g2_decap_8
XFILLER_20_497 VDD VSS sg13g2_decap_8
XFILLER_106_525 VDD VSS sg13g2_decap_8
XFILLER_109_7 VDD VSS sg13g2_decap_8
XFILLER_88_921 VDD VSS sg13g2_decap_8
XFILLER_102_731 VDD VSS sg13g2_fill_1
XFILLER_0_847 VDD VSS sg13g2_decap_8
XFILLER_58_14 VDD VSS sg13g2_decap_8
XFILLER_88_965 VDD VSS sg13g2_decap_8
XFILLER_101_241 VDD VSS sg13g2_decap_8
XFILLER_48_807 VDD VSS sg13g2_decap_8
XFILLER_75_637 VDD VSS sg13g2_decap_8
XFILLER_87_475 VDD VSS sg13g2_decap_8
XFILLER_74_147 VDD VSS sg13g2_decap_8
XFILLER_90_629 VDD VSS sg13g2_fill_1
XFILLER_83_670 VDD VSS sg13g2_decap_8
XFILLER_74_35 VDD VSS sg13g2_decap_8
XFILLER_28_553 VDD VSS sg13g2_decap_8
XFILLER_62_309 VDD VSS sg13g2_decap_8
XFILLER_55_361 VDD VSS sg13g2_decap_8
XFILLER_70_320 VDD VSS sg13g2_decap_8
XFILLER_55_372 VDD VSS sg13g2_fill_2
XFILLER_15_203 VDD VSS sg13g2_decap_8
XFILLER_43_512 VDD VSS sg13g2_decap_4
XFILLER_71_854 VDD VSS sg13g2_decap_8
XFILLER_43_545 VDD VSS sg13g2_decap_8
XFILLER_31_707 VDD VSS sg13g2_decap_8
XFILLER_70_386 VDD VSS sg13g2_decap_8
XFILLER_24_770 VDD VSS sg13g2_decap_8
XFILLER_12_910 VDD VSS sg13g2_decap_8
XFILLER_30_217 VDD VSS sg13g2_decap_8
XFILLER_90_56 VDD VSS sg13g2_decap_8
XFILLER_11_420 VDD VSS sg13g2_decap_8
XFILLER_8_903 VDD VSS sg13g2_decap_8
XFILLER_23_280 VDD VSS sg13g2_decap_8
XFILLER_7_413 VDD VSS sg13g2_decap_8
XFILLER_12_987 VDD VSS sg13g2_decap_8
XFILLER_99_21 VDD VSS sg13g2_decap_8
XFILLER_11_497 VDD VSS sg13g2_decap_8
XFILLER_87_1054 VDD VSS sg13g2_decap_8
XFILLER_99_98 VDD VSS sg13g2_decap_8
XFILLER_48_1016 VDD VSS sg13g2_decap_8
XFILLER_3_630 VDD VSS sg13g2_decap_8
XFILLER_98_718 VDD VSS sg13g2_decap_8
X_2363__281 VDD VSS _2363_/RESET_B sg13g2_tiehi
XFILLER_2_140 VDD VSS sg13g2_decap_8
XFILLER_112_539 VDD VSS sg13g2_decap_8
XFILLER_97_228 VDD VSS sg13g2_decap_8
XFILLER_79_954 VDD VSS sg13g2_decap_8
XFILLER_94_913 VDD VSS sg13g2_decap_8
XFILLER_24_7 VDD VSS sg13g2_decap_8
XFILLER_66_637 VDD VSS sg13g2_fill_2
XFILLER_39_829 VDD VSS sg13g2_decap_8
XFILLER_38_306 VDD VSS sg13g2_decap_8
XFILLER_93_456 VDD VSS sg13g2_decap_8
X_2090_ _2149_/B _2082_/B _2085_/X _2343_/D VDD VSS sg13g2_a21o_1
XFILLER_81_629 VDD VSS sg13g2_decap_8
XFILLER_47_873 VDD VSS sg13g2_decap_8
XFILLER_47_884 VDD VSS sg13g2_fill_1
XFILLER_0_21 VDD VSS sg13g2_decap_8
XFILLER_19_553 VDD VSS sg13g2_decap_8
XFILLER_94_1025 VDD VSS sg13g2_decap_4
XFILLER_74_681 VDD VSS sg13g2_decap_8
XFILLER_62_843 VDD VSS sg13g2_decap_8
XFILLER_0_1029 VDD VSS sg13g2_decap_8
XFILLER_34_567 VDD VSS sg13g2_decap_8
XFILLER_22_707 VDD VSS sg13g2_decap_8
XFILLER_0_98 VDD VSS sg13g2_decap_8
XFILLER_15_770 VDD VSS sg13g2_decap_8
XFILLER_21_217 VDD VSS sg13g2_decap_8
X_1943_ _1946_/A _1943_/A _1943_/B VDD VSS sg13g2_xnor2_1
XFILLER_61_397 VDD VSS sg13g2_decap_8
XFILLER_14_280 VDD VSS sg13g2_decap_8
XFILLER_9_63 VDD VSS sg13g2_decap_8
XFILLER_30_784 VDD VSS sg13g2_decap_8
X_1874_ _1884_/B _1874_/A _1874_/B VDD VSS sg13g2_xnor2_1
XIO_FILL_IO_SOUTH_5_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_2288__157 VDD VSS _2288_/RESET_B sg13g2_tiehi
XFILLER_7_980 VDD VSS sg13g2_decap_8
XFILLER_6_490 VDD VSS sg13g2_decap_8
XFILLER_50_0 VDD VSS sg13g2_decap_8
XFILLER_103_517 VDD VSS sg13g2_decap_8
XFILLER_88_206 VDD VSS sg13g2_decap_8
XFILLER_69_431 VDD VSS sg13g2_fill_1
XFILLER_9_1043 VDD VSS sg13g2_decap_8
XFILLER_57_604 VDD VSS sg13g2_decap_8
XFILLER_28_28 VDD VSS sg13g2_decap_8
XFILLER_56_103 VDD VSS sg13g2_decap_8
X_2357_ _2357_/RESET_B VSS VDD _2357_/D _2357_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_85_957 VDD VSS sg13g2_decap_8
X_1308_ _1308_/Y _1342_/B1 hold385/X _1342_/A2 _2348_/Q VDD VSS sg13g2_a22oi_1
XFILLER_96_294 VDD VSS sg13g2_decap_8
X_2288_ _2288_/RESET_B VSS VDD _2288_/D _2288_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_84_489 VDD VSS sg13g2_decap_8
XFILLER_53_810 VDD VSS sg13g2_decap_8
XFILLER_38_884 VDD VSS sg13g2_decap_8
X_1239_ _1248_/A _2297_/Q _2259_/Q VDD VSS sg13g2_xnor2_1
XFILLER_37_350 VDD VSS sg13g2_decap_8
XFILLER_25_567 VDD VSS sg13g2_decap_8
XFILLER_13_707 VDD VSS sg13g2_decap_8
XFILLER_44_49 VDD VSS sg13g2_decap_8
X_2236__270 VDD VSS _2236_/RESET_B sg13g2_tiehi
XFILLER_53_898 VDD VSS sg13g2_fill_2
XFILLER_53_887 VDD VSS sg13g2_decap_8
XFILLER_52_375 VDD VSS sg13g2_decap_8
XFILLER_12_217 VDD VSS sg13g2_decap_8
XFILLER_40_526 VDD VSS sg13g2_decap_4
XFILLER_40_537 VDD VSS sg13g2_fill_1
XFILLER_100_77 VDD VSS sg13g2_decap_8
XFILLER_21_784 VDD VSS sg13g2_decap_8
XFILLER_60_59 VDD VSS sg13g2_decap_8
X_2267__219 VDD VSS _2267_/RESET_B sg13g2_tiehi
XFILLER_20_294 VDD VSS sg13g2_decap_8
XFILLER_5_917 VDD VSS sg13g2_decap_8
XFILLER_107_856 VDD VSS sg13g2_decap_8
XFILLER_106_333 VDD VSS sg13g2_decap_8
XFILLER_109_42 VDD VSS sg13g2_decap_8
XFILLER_4_427 VDD VSS sg13g2_decap_8
XFILLER_106_344 VDD VSS sg13g2_fill_2
XFILLER_69_35 VDD VSS sg13g2_decap_8
XFILLER_79_217 VDD VSS sg13g2_decap_8
XFILLER_0_644 VDD VSS sg13g2_decap_8
XFILLER_88_795 VDD VSS sg13g2_decap_8
XFILLER_87_283 VDD VSS sg13g2_decap_8
XFILLER_85_56 VDD VSS sg13g2_decap_8
XFILLER_48_659 VDD VSS sg13g2_decap_8
XFILLER_29_840 VDD VSS sg13g2_decap_8
XFILLER_47_125 VDD VSS sg13g2_decap_8
XFILLER_63_607 VDD VSS sg13g2_decap_8
XFILLER_28_350 VDD VSS sg13g2_decap_8
XFILLER_44_832 VDD VSS sg13g2_decap_4
XFILLER_71_640 VDD VSS sg13g2_decap_8
XFILLER_44_865 VDD VSS sg13g2_decap_8
XFILLER_16_567 VDD VSS sg13g2_decap_8
XFILLER_71_684 VDD VSS sg13g2_fill_1
XFILLER_70_161 VDD VSS sg13g2_decap_8
XFILLER_31_504 VDD VSS sg13g2_decap_8
XFILLER_43_364 VDD VSS sg13g2_decap_8
XFILLER_8_700 VDD VSS sg13g2_decap_8
XFILLER_15_1015 VDD VSS sg13g2_decap_8
XFILLER_7_210 VDD VSS sg13g2_decap_8
XFILLER_12_784 VDD VSS sg13g2_decap_8
XFILLER_11_294 VDD VSS sg13g2_decap_8
XFILLER_8_777 VDD VSS sg13g2_decap_8
XFILLER_109_182 VDD VSS sg13g2_fill_2
XFILLER_7_287 VDD VSS sg13g2_decap_8
XFILLER_50_92 VDD VSS sg13g2_decap_8
X_1590_ _1595_/A _1590_/B _1592_/B _2287_/D VDD VSS sg13g2_nor3_1
XFILLER_98_504 VDD VSS sg13g2_decap_8
XFILLER_4_994 VDD VSS sg13g2_decap_8
XFILLER_112_336 VDD VSS sg13g2_decap_8
X_2211_ _2211_/RESET_B VSS VDD _2211_/D _2211_/Q clkload5/A sg13g2_dfrbpq_1
XFILLER_39_626 VDD VSS sg13g2_decap_8
X_2142_ _2071_/A VDD _2143_/B VSS _2142_/A1 hold565/X sg13g2_o21ai_1
XFILLER_93_220 VDD VSS sg13g2_fill_1
XFILLER_67_957 VDD VSS sg13g2_decap_8
XFILLER_22_1008 VDD VSS sg13g2_decap_8
X_2073_ _2063_/X _2086_/A _2079_/S _2074_/B VDD VSS sg13g2_mux2_1
XFILLER_93_264 VDD VSS sg13g2_fill_2
XFILLER_66_456 VDD VSS sg13g2_decap_8
XFILLER_19_350 VDD VSS sg13g2_decap_8
XFILLER_38_147 VDD VSS sg13g2_decap_8
XFILLER_82_949 VDD VSS sg13g2_decap_8
XFILLER_81_426 VDD VSS sg13g2_decap_8
XFILLER_53_139 VDD VSS sg13g2_decap_8
XFILLER_35_854 VDD VSS sg13g2_decap_8
XFILLER_62_662 VDD VSS sg13g2_decap_8
XFILLER_61_150 VDD VSS sg13g2_decap_8
XFILLER_22_504 VDD VSS sg13g2_decap_8
XFILLER_34_364 VDD VSS sg13g2_decap_8
XFILLER_98_0 VDD VSS sg13g2_decap_8
XFILLER_50_857 VDD VSS sg13g2_decap_4
X_1926_ _1928_/A _1926_/A _1926_/B VDD VSS sg13g2_xnor2_1
XFILLER_30_581 VDD VSS sg13g2_decap_8
X_1857_ _2003_/A _2244_/Q _2203_/Q VDD VSS sg13g2_xnor2_1
XFILLER_107_119 VDD VSS sg13g2_decap_8
Xfanout4 _2074_/A _2149_/A VDD VSS sg13g2_buf_1
X_1788_ _1900_/B _1912_/B _1817_/B VDD VSS sg13g2_and2_1
XFILLER_89_537 VDD VSS sg13g2_decap_8
XFILLER_89_515 VDD VSS sg13g2_decap_8
XFILLER_97_570 VDD VSS sg13g2_decap_8
XFILLER_85_721 VDD VSS sg13g2_decap_8
XFILLER_103_369 VDD VSS sg13g2_decap_8
XFILLER_39_49 VDD VSS sg13g2_decap_8
XFILLER_58_957 VDD VSS sg13g2_fill_2
XFILLER_84_264 VDD VSS sg13g2_decap_8
XFILLER_29_147 VDD VSS sg13g2_decap_8
XFILLER_85_798 VDD VSS sg13g2_decap_8
XFILLER_38_681 VDD VSS sg13g2_decap_8
XFILLER_81_960 VDD VSS sg13g2_decap_8
XFILLER_77_1042 VDD VSS sg13g2_decap_8
XFILLER_111_21 VDD VSS sg13g2_decap_8
XFILLER_26_854 VDD VSS sg13g2_decap_8
XFILLER_53_673 VDD VSS sg13g2_decap_4
XFILLER_13_504 VDD VSS sg13g2_decap_8
XFILLER_25_364 VDD VSS sg13g2_decap_8
XFILLER_80_481 VDD VSS sg13g2_decap_8
XFILLER_111_98 VDD VSS sg13g2_decap_8
XFILLER_71_14 VDD VSS sg13g2_decap_8
XFILLER_38_1059 VDD VSS sg13g2_fill_2
XFILLER_41_846 VDD VSS sg13g2_decap_8
XFILLER_40_356 VDD VSS sg13g2_decap_8
XFILLER_21_581 VDD VSS sg13g2_decap_8
XFILLER_5_714 VDD VSS sg13g2_decap_8
XFILLER_4_224 VDD VSS sg13g2_decap_8
XFILLER_107_653 VDD VSS sg13g2_decap_8
XFILLER_20_84 VDD VSS sg13g2_decap_8
XFILLER_106_196 VDD VSS sg13g2_decap_8
XFILLER_1_931 VDD VSS sg13g2_decap_8
XIO_BOND_in_data_pads\[6\].in_data_pad in_data_PADs[6] bondpad_70x70
XFILLER_103_870 VDD VSS sg13g2_fill_1
X_2321__224 VDD VSS _2321_/RESET_B sg13g2_tiehi
XFILLER_95_529 VDD VSS sg13g2_decap_8
XFILLER_96_77 VDD VSS sg13g2_decap_8
XFILLER_49_924 VDD VSS sg13g2_decap_8
XFILLER_67_209 VDD VSS sg13g2_decap_8
XFILLER_0_441 VDD VSS sg13g2_decap_8
XFILLER_48_423 VDD VSS sg13g2_decap_8
XFILLER_76_776 VDD VSS sg13g2_decap_8
XFILLER_75_264 VDD VSS sg13g2_decap_8
XFILLER_63_415 VDD VSS sg13g2_decap_4
XFILLER_63_426 VDD VSS sg13g2_decap_8
XFILLER_48_489 VDD VSS sg13g2_decap_8
XFILLER_90_256 VDD VSS sg13g2_decap_8
XFILLER_17_854 VDD VSS sg13g2_decap_8
XFILLER_16_364 VDD VSS sg13g2_decap_8
XFILLER_45_70 VDD VSS sg13g2_decap_8
XFILLER_31_301 VDD VSS sg13g2_decap_8
XFILLER_91_1028 VDD VSS sg13g2_decap_8
XFILLER_71_481 VDD VSS sg13g2_decap_8
XFILLER_91_7 VDD VSS sg13g2_decap_8
XFILLER_32_868 VDD VSS sg13g2_decap_8
XFILLER_31_378 VDD VSS sg13g2_decap_8
XFILLER_12_581 VDD VSS sg13g2_decap_8
X_1711_ _1710_/Y VDD _1711_/Y VSS _1720_/A hold514/X sg13g2_o21ai_1
XFILLER_8_574 VDD VSS sg13g2_decap_8
X_1642_ _1671_/D _1677_/A _1674_/B VDD VSS sg13g2_nand2_1
XFILLER_6_42 VDD VSS sg13g2_decap_8
X_1573_ _1572_/Y VDD _1573_/Y VSS _1573_/A1 _2209_/Q sg13g2_o21ai_1
XFILLER_101_807 VDD VSS sg13g2_decap_8
XFILLER_99_857 VDD VSS sg13g2_decap_8
XFILLER_112_133 VDD VSS sg13g2_decap_8
XFILLER_4_791 VDD VSS sg13g2_decap_8
XFILLER_98_367 VDD VSS sg13g2_fill_1
XFILLER_39_401 VDD VSS sg13g2_decap_8
XFILLER_82_702 VDD VSS sg13g2_decap_8
XFILLER_55_916 VDD VSS sg13g2_decap_4
XFILLER_67_776 VDD VSS sg13g2_decap_8
XFILLER_13_0 VDD VSS sg13g2_decap_8
XFILLER_6_1057 VDD VSS sg13g2_decap_4
XFILLER_39_478 VDD VSS sg13g2_decap_8
X_2125_ VDD VSS hold325/X _2120_/A _2124_/Y _2124_/B _2127_/A _2123_/X sg13g2_a221oi_1
XFILLER_94_573 VDD VSS sg13g2_decap_8
XFILLER_66_264 VDD VSS sg13g2_decap_8
XFILLER_54_404 VDD VSS sg13g2_decap_8
X_2056_ _1908_/A _1922_/Y _2069_/S _2056_/X VDD VSS sg13g2_mux2_1
XFILLER_81_256 VDD VSS sg13g2_decap_8
XFILLER_35_651 VDD VSS sg13g2_decap_8
XFILLER_62_470 VDD VSS sg13g2_decap_8
XFILLER_34_161 VDD VSS sg13g2_decap_8
XFILLER_22_301 VDD VSS sg13g2_decap_8
XFILLER_50_643 VDD VSS sg13g2_decap_8
XFILLER_23_868 VDD VSS sg13g2_decap_8
XFILLER_10_518 VDD VSS sg13g2_decap_8
XFILLER_41_28 VDD VSS sg13g2_decap_8
XFILLER_22_378 VDD VSS sg13g2_decap_8
X_1909_ _1907_/B _1908_/Y _1954_/S _1943_/B VDD VSS sg13g2_mux2_1
Xhold530 _2271_/Q VDD VSS hold530/X sg13g2_dlygate4sd3_1
Xhold541 _1718_/Y VDD VSS _2318_/D sg13g2_dlygate4sd3_1
XFILLER_104_612 VDD VSS sg13g2_decap_8
XFILLER_2_728 VDD VSS sg13g2_decap_8
Xhold563 _1639_/Y VDD VSS _2297_/D sg13g2_dlygate4sd3_1
Xhold552 _1620_/Y VDD VSS _1621_/B sg13g2_dlygate4sd3_1
XFILLER_89_356 VDD VSS sg13g2_decap_8
XFILLER_103_133 VDD VSS sg13g2_decap_8
XFILLER_1_238 VDD VSS sg13g2_decap_8
XFILLER_104_689 VDD VSS sg13g2_decap_8
XFILLER_89_367 VDD VSS sg13g2_fill_1
XFILLER_106_21 VDD VSS sg13g2_decap_8
XFILLER_58_721 VDD VSS sg13g2_decap_8
XFILLER_66_14 VDD VSS sg13g2_decap_8
XFILLER_100_840 VDD VSS sg13g2_decap_8
XFILLER_85_540 VDD VSS sg13g2_decap_8
XFILLER_106_98 VDD VSS sg13g2_decap_8
XFILLER_57_253 VDD VSS sg13g2_decap_4
XFILLER_39_990 VDD VSS sg13g2_decap_8
XFILLER_57_297 VDD VSS sg13g2_decap_8
XFILLER_45_448 VDD VSS sg13g2_decap_8
XFILLER_45_437 VDD VSS sg13g2_fill_2
XFILLER_82_35 VDD VSS sg13g2_decap_8
XFILLER_26_651 VDD VSS sg13g2_decap_8
XFILLER_60_429 VDD VSS sg13g2_decap_8
XFILLER_41_643 VDD VSS sg13g2_decap_8
XFILLER_53_470 VDD VSS sg13g2_decap_8
XFILLER_13_301 VDD VSS sg13g2_decap_8
XFILLER_25_161 VDD VSS sg13g2_decap_8
XFILLER_15_84 VDD VSS sg13g2_decap_8
XFILLER_14_868 VDD VSS sg13g2_decap_8
XFILLER_90_1050 VDD VSS sg13g2_decap_8
XFILLER_13_378 VDD VSS sg13g2_decap_8
XFILLER_40_175 VDD VSS sg13g2_decap_8
XFILLER_51_1045 VDD VSS sg13g2_decap_8
XFILLER_5_511 VDD VSS sg13g2_decap_8
XFILLER_12_1029 VDD VSS sg13g2_decap_8
XFILLER_108_962 VDD VSS sg13g2_decap_8
Xiovdd_pads\[0\].iovdd_pad IOVDD IOVSS VDD VSS sg13g2_IOPadIOVdd
XFILLER_107_472 VDD VSS sg13g2_decap_8
XFILLER_107_483 VDD VSS sg13g2_fill_1
XFILLER_5_588 VDD VSS sg13g2_decap_8
XFILLER_107_494 VDD VSS sg13g2_fill_2
X_2206__128 VDD VSS _2206_/RESET_B sg13g2_tiehi
XFILLER_110_648 VDD VSS sg13g2_decap_8
X_2180__180 VDD VSS _2180_/RESET_B sg13g2_tiehi
XFILLER_76_540 VDD VSS sg13g2_decap_8
XFILLER_49_776 VDD VSS sg13g2_decap_8
XFILLER_48_253 VDD VSS sg13g2_decap_8
XFILLER_91_521 VDD VSS sg13g2_decap_8
XFILLER_37_938 VDD VSS sg13g2_decap_8
XFILLER_64_746 VDD VSS sg13g2_decap_8
XFILLER_52_908 VDD VSS sg13g2_decap_8
XFILLER_36_448 VDD VSS sg13g2_decap_8
XFILLER_45_982 VDD VSS sg13g2_decap_8
XFILLER_51_429 VDD VSS sg13g2_decap_8
XFILLER_17_651 VDD VSS sg13g2_decap_8
XFILLER_91_598 VDD VSS sg13g2_fill_1
XFILLER_16_161 VDD VSS sg13g2_decap_8
XFILLER_44_481 VDD VSS sg13g2_decap_8
XFILLER_108_1046 VDD VSS sg13g2_decap_8
XFILLER_60_963 VDD VSS sg13g2_decap_8
XFILLER_32_665 VDD VSS sg13g2_decap_8
XFILLER_20_805 VDD VSS sg13g2_decap_8
XFILLER_31_175 VDD VSS sg13g2_decap_8
XFILLER_9_861 VDD VSS sg13g2_decap_8
XFILLER_8_371 VDD VSS sg13g2_decap_8
X_1625_ _1624_/Y VDD _1625_/Y VSS _1634_/A hold500/X sg13g2_o21ai_1
XFILLER_99_632 VDD VSS sg13g2_decap_8
X_1556_ _1556_/S0 _2239_/Q _2231_/Q _2223_/Q _2215_/Q _1589_/B _1557_/A VDD VSS sg13g2_mux4_1
XFILLER_101_615 VDD VSS sg13g2_decap_8
XFILLER_99_687 VDD VSS sg13g2_decap_8
XFILLER_28_1036 VDD VSS sg13g2_decap_8
XFILLER_59_518 VDD VSS sg13g2_decap_8
XFILLER_101_648 VDD VSS sg13g2_decap_8
XFILLER_98_197 VDD VSS sg13g2_decap_8
X_1487_ _1487_/Y _1487_/A _1487_/B VDD VSS sg13g2_nand2_1
XFILLER_100_147 VDD VSS sg13g2_decap_8
XFILLER_39_231 VDD VSS sg13g2_fill_2
XFILLER_95_882 VDD VSS sg13g2_decap_8
XFILLER_28_938 VDD VSS sg13g2_decap_8
XFILLER_67_595 VDD VSS sg13g2_decap_8
XFILLER_55_713 VDD VSS sg13g2_decap_8
XFILLER_36_28 VDD VSS sg13g2_decap_8
XFILLER_54_245 VDD VSS sg13g2_decap_8
XFILLER_27_448 VDD VSS sg13g2_decap_8
X_2108_ VSS VDD _1220_/A _2106_/B _2108_/Y _2107_/Y sg13g2_a21oi_1
XFILLER_82_576 VDD VSS sg13g2_decap_8
XFILLER_43_919 VDD VSS sg13g2_decap_8
XFILLER_54_256 VDD VSS sg13g2_fill_2
X_2039_ _2038_/X _2082_/B _2037_/X _2326_/D VDD VSS sg13g2_a21o_1
XFILLER_70_738 VDD VSS sg13g2_decap_8
XFILLER_74_1045 VDD VSS sg13g2_decap_8
XFILLER_35_1029 VDD VSS sg13g2_decap_8
XFILLER_23_665 VDD VSS sg13g2_decap_8
XFILLER_11_805 VDD VSS sg13g2_decap_8
XFILLER_50_451 VDD VSS sg13g2_decap_8
XFILLER_51_996 VDD VSS sg13g2_decap_8
XFILLER_10_315 VDD VSS sg13g2_decap_8
XFILLER_22_175 VDD VSS sg13g2_decap_8
XFILLER_6_308 VDD VSS sg13g2_decap_8
XFILLER_108_214 VDD VSS sg13g2_decap_4
XFILLER_108_236 VDD VSS sg13g2_decap_8
XFILLER_105_910 VDD VSS sg13g2_decap_8
Xhold360 _2175_/Q VDD VSS hold360/X sg13g2_dlygate4sd3_1
Xhold371 _2309_/Q VDD VSS _1225_/B sg13g2_dlygate4sd3_1
XFILLER_2_525 VDD VSS sg13g2_decap_8
XFILLER_105_987 VDD VSS sg13g2_decap_8
XFILLER_78_827 VDD VSS sg13g2_decap_8
Xhold382 _1328_/Y VDD VSS _1329_/A sg13g2_dlygate4sd3_1
XFILLER_77_35 VDD VSS sg13g2_decap_8
Xhold393 _1486_/Y VDD VSS _2263_/D sg13g2_dlygate4sd3_1
XFILLER_89_186 VDD VSS sg13g2_decap_8
XFILLER_77_315 VDD VSS sg13g2_decap_8
XFILLER_19_938 VDD VSS sg13g2_decap_8
XFILLER_93_56 VDD VSS sg13g2_decap_8
XFILLER_46_768 VDD VSS sg13g2_decap_8
XFILLER_18_448 VDD VSS sg13g2_decap_8
XFILLER_42_952 VDD VSS sg13g2_decap_8
XFILLER_14_665 VDD VSS sg13g2_decap_8
XFILLER_41_451 VDD VSS sg13g2_decap_8
XFILLER_13_175 VDD VSS sg13g2_decap_8
XFILLER_41_495 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_6_2 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_9_168 VDD VSS sg13g2_decap_8
XFILLER_10_882 VDD VSS sg13g2_decap_8
XFILLER_6_875 VDD VSS sg13g2_decap_8
XFILLER_54_7 VDD VSS sg13g2_decap_8
XFILLER_107_291 VDD VSS sg13g2_decap_8
X_1410_ _1410_/Y _2265_/Q _1410_/B VDD VSS sg13g2_nand2_1
XFILLER_5_385 VDD VSS sg13g2_decap_8
XFILLER_69_816 VDD VSS sg13g2_decap_8
Xvdd_pads\[0\].vdd_pad IOVDD IOVSS VDD VSS sg13g2_IOPadVdd
XFILLER_3_21 VDD VSS sg13g2_decap_8
XFILLER_111_924 VDD VSS sg13g2_decap_8
X_1341_ VDD _2200_/D _1341_/A VSS sg13g2_inv_1
XFILLER_95_112 VDD VSS sg13g2_decap_8
XFILLER_68_326 VDD VSS sg13g2_decap_8
X_1272_ _1272_/Y _1338_/B1 hold345/X _1338_/A2 _2316_/Q VDD VSS sg13g2_a22oi_1
XFILLER_96_679 VDD VSS sg13g2_decap_8
XFILLER_110_445 VDD VSS sg13g2_decap_8
XFILLER_49_551 VDD VSS sg13g2_decap_8
XFILLER_3_98 VDD VSS sg13g2_decap_8
XFILLER_95_189 VDD VSS sg13g2_decap_8
XFILLER_64_543 VDD VSS sg13g2_decap_8
XFILLER_37_735 VDD VSS sg13g2_decap_8
XFILLER_91_362 VDD VSS sg13g2_fill_2
XFILLER_52_705 VDD VSS sg13g2_decap_8
XFILLER_36_245 VDD VSS sg13g2_decap_8
XIO_FILL_IO_NORTH_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_52_738 VDD VSS sg13g2_fill_1
XFILLER_45_790 VDD VSS sg13g2_decap_4
XFILLER_51_237 VDD VSS sg13g2_decap_8
XFILLER_33_952 VDD VSS sg13g2_decap_8
XFILLER_60_771 VDD VSS sg13g2_decap_8
XFILLER_20_602 VDD VSS sg13g2_decap_8
XFILLER_32_462 VDD VSS sg13g2_decap_8
XFILLER_80_0 VDD VSS sg13g2_decap_8
XFILLER_20_679 VDD VSS sg13g2_decap_8
XFILLER_105_228 VDD VSS sg13g2_decap_8
X_1608_ _1608_/Y _1638_/S _1612_/A VDD VSS sg13g2_nand2_1
XFILLER_102_902 VDD VSS sg13g2_decap_8
XFILLER_99_462 VDD VSS sg13g2_decap_8
XFILLER_102_935 VDD VSS sg13g2_decap_8
XFILLER_101_423 VDD VSS sg13g2_decap_8
X_1539_ _1538_/Y VDD _1539_/Y VSS _1592_/A _1536_/Y sg13g2_o21ai_1
XFILLER_87_668 VDD VSS sg13g2_decap_8
XFILLER_41_1000 VDD VSS sg13g2_decap_8
XFILLER_59_348 VDD VSS sg13g2_decap_8
XFILLER_86_178 VDD VSS sg13g2_decap_8
XFILLER_74_307 VDD VSS sg13g2_decap_8
XFILLER_47_49 VDD VSS sg13g2_decap_8
XFILLER_83_841 VDD VSS sg13g2_decap_4
XFILLER_28_735 VDD VSS sg13g2_decap_8
XFILLER_67_381 VDD VSS sg13g2_decap_4
XFILLER_83_885 VDD VSS sg13g2_decap_8
XFILLER_43_716 VDD VSS sg13g2_decap_8
XFILLER_27_245 VDD VSS sg13g2_decap_8
XFILLER_70_535 VDD VSS sg13g2_decap_8
XFILLER_103_77 VDD VSS sg13g2_decap_8
XFILLER_42_226 VDD VSS sg13g2_fill_1
XFILLER_24_952 VDD VSS sg13g2_decap_8
XFILLER_42_259 VDD VSS sg13g2_decap_8
XFILLER_51_793 VDD VSS sg13g2_decap_8
XFILLER_11_602 VDD VSS sg13g2_decap_8
XFILLER_23_462 VDD VSS sg13g2_decap_8
XFILLER_10_112 VDD VSS sg13g2_decap_8
XFILLER_6_105 VDD VSS sg13g2_decap_8
XFILLER_11_679 VDD VSS sg13g2_decap_8
XFILLER_109_567 VDD VSS sg13g2_decap_8
XFILLER_10_189 VDD VSS sg13g2_decap_8
XFILLER_12_63 VDD VSS sg13g2_decap_8
XFILLER_3_812 VDD VSS sg13g2_decap_8
XFILLER_2_322 VDD VSS sg13g2_decap_8
XFILLER_78_602 VDD VSS sg13g2_decap_8
XFILLER_88_56 VDD VSS sg13g2_decap_8
XFILLER_3_889 VDD VSS sg13g2_decap_8
XFILLER_105_784 VDD VSS sg13g2_decap_8
XFILLER_78_635 VDD VSS sg13g2_fill_1
XFILLER_77_112 VDD VSS sg13g2_decap_8
XFILLER_2_399 VDD VSS sg13g2_decap_8
XFILLER_77_189 VDD VSS sg13g2_decap_8
X_2306__87 VDD VSS _2306__87/L_HI sg13g2_tiehi
XFILLER_65_329 VDD VSS sg13g2_fill_1
XFILLER_46_510 VDD VSS sg13g2_decap_8
XFILLER_93_649 VDD VSS sg13g2_decap_8
XFILLER_58_392 VDD VSS sg13g2_decap_8
XFILLER_19_735 VDD VSS sg13g2_decap_8
XFILLER_74_863 VDD VSS sg13g2_fill_2
XFILLER_73_351 VDD VSS sg13g2_decap_8
XFILLER_18_245 VDD VSS sg13g2_decap_8
XFILLER_34_749 VDD VSS sg13g2_decap_8
XFILLER_61_557 VDD VSS sg13g2_decap_4
XFILLER_15_952 VDD VSS sg13g2_decap_8
XFILLER_33_259 VDD VSS sg13g2_decap_8
XFILLER_14_462 VDD VSS sg13g2_decap_8
X_1890_ _1895_/A _1891_/A _1891_/B VDD VSS sg13g2_nand2_1
XFILLER_30_966 VDD VSS sg13g2_decap_8
XFILLER_18_1057 VDD VSS sg13g2_decap_4
XFILLER_41_281 VDD VSS sg13g2_fill_2
XFILLER_6_672 VDD VSS sg13g2_decap_8
XFILLER_5_182 VDD VSS sg13g2_decap_8
XFILLER_102_209 VDD VSS sg13g2_fill_1
XFILLER_64_1000 VDD VSS sg13g2_decap_8
XFILLER_97_944 VDD VSS sg13g2_decap_4
XFILLER_111_721 VDD VSS sg13g2_decap_8
XFILLER_69_635 VDD VSS sg13g2_decap_8
X_2373_ _2373__93/L_HI VSS VDD _2373_/D _2373_/Q _2373_/CLK sg13g2_dfrbpq_1
XFILLER_97_977 VDD VSS sg13g2_decap_8
X_1324_ _1324_/Y _1342_/B1 hold343/X _1342_/A2 _2325_/Q VDD VSS sg13g2_a22oi_1
XFILLER_110_231 VDD VSS sg13g2_decap_8
XFILLER_111_798 VDD VSS sg13g2_decap_8
XFILLER_84_627 VDD VSS sg13g2_decap_8
XFILLER_83_137 VDD VSS sg13g2_fill_1
XFILLER_83_126 VDD VSS sg13g2_decap_8
XFILLER_65_841 VDD VSS sg13g2_decap_4
X_1255_ _1260_/A _1255_/B _1507_/A VDD VSS sg13g2_nor2_1
XFILLER_37_532 VDD VSS sg13g2_decap_8
XFILLER_92_682 VDD VSS sg13g2_decap_8
XFILLER_25_749 VDD VSS sg13g2_decap_8
XFILLER_64_395 VDD VSS sg13g2_decap_8
XFILLER_91_192 VDD VSS sg13g2_decap_8
XFILLER_24_259 VDD VSS sg13g2_decap_8
XFILLER_71_1026 VDD VSS sg13g2_decap_8
XFILLER_21_966 VDD VSS sg13g2_decap_8
XFILLER_60_590 VDD VSS sg13g2_decap_4
XFILLER_20_476 VDD VSS sg13g2_decap_8
XFILLER_106_504 VDD VSS sg13g2_decap_8
XFILLER_4_609 VDD VSS sg13g2_decap_8
XFILLER_3_119 VDD VSS sg13g2_decap_8
XFILLER_106_559 VDD VSS sg13g2_decap_8
XFILLER_88_900 VDD VSS sg13g2_decap_8
XFILLER_99_270 VDD VSS sg13g2_decap_4
XFILLER_0_826 VDD VSS sg13g2_decap_8
XFILLER_101_220 VDD VSS sg13g2_decap_8
XFILLER_59_145 VDD VSS sg13g2_fill_2
XFILLER_102_787 VDD VSS sg13g2_fill_2
XFILLER_75_616 VDD VSS sg13g2_decap_8
XFILLER_101_297 VDD VSS sg13g2_fill_1
XFILLER_74_126 VDD VSS sg13g2_decap_8
XFILLER_74_14 VDD VSS sg13g2_decap_8
XFILLER_28_532 VDD VSS sg13g2_decap_8
XFILLER_90_608 VDD VSS sg13g2_decap_8
XFILLER_56_885 VDD VSS sg13g2_decap_8
XFILLER_71_833 VDD VSS sg13g2_decap_8
XFILLER_82_170 VDD VSS sg13g2_fill_2
XFILLER_16_749 VDD VSS sg13g2_decap_8
XFILLER_43_535 VDD VSS sg13g2_decap_4
XFILLER_15_259 VDD VSS sg13g2_decap_8
XFILLER_70_365 VDD VSS sg13g2_decap_8
XFILLER_90_35 VDD VSS sg13g2_decap_8
XFILLER_12_966 VDD VSS sg13g2_decap_8
XFILLER_109_320 VDD VSS sg13g2_decap_4
XFILLER_11_476 VDD VSS sg13g2_decap_8
XFILLER_8_959 VDD VSS sg13g2_decap_8
XFILLER_23_84 VDD VSS sg13g2_decap_8
XFILLER_7_469 VDD VSS sg13g2_decap_8
XFILLER_99_77 VDD VSS sg13g2_decap_8
XFILLER_97_207 VDD VSS sg13g2_decap_8
XFILLER_105_581 VDD VSS sg13g2_decap_8
XFILLER_112_518 VDD VSS sg13g2_decap_8
XFILLER_78_410 VDD VSS sg13g2_decap_8
XFILLER_3_686 VDD VSS sg13g2_decap_8
XFILLER_78_443 VDD VSS sg13g2_decap_8
XFILLER_78_454 VDD VSS sg13g2_fill_2
XFILLER_39_808 VDD VSS sg13g2_decap_8
XFILLER_2_196 VDD VSS sg13g2_decap_8
XFILLER_66_616 VDD VSS sg13g2_decap_8
XFILLER_94_969 VDD VSS sg13g2_decap_8
XFILLER_93_435 VDD VSS sg13g2_decap_8
XFILLER_24_1050 VDD VSS sg13g2_decap_8
XFILLER_17_7 VDD VSS sg13g2_decap_8
XFILLER_19_532 VDD VSS sg13g2_decap_8
XFILLER_81_608 VDD VSS sg13g2_decap_8
XFILLER_74_660 VDD VSS sg13g2_decap_8
XFILLER_0_1008 VDD VSS sg13g2_decap_8
XFILLER_65_148 VDD VSS sg13g2_fill_2
XFILLER_46_340 VDD VSS sg13g2_decap_8
XFILLER_94_1004 VDD VSS sg13g2_decap_8
XFILLER_62_822 VDD VSS sg13g2_decap_8
XFILLER_0_77 VDD VSS sg13g2_decap_8
XFILLER_94_1059 VDD VSS sg13g2_fill_2
XFILLER_94_1048 VDD VSS sg13g2_decap_8
XFILLER_34_546 VDD VSS sg13g2_decap_8
XFILLER_61_354 VDD VSS sg13g2_decap_8
XFILLER_62_899 VDD VSS sg13g2_decap_8
X_1942_ _1992_/B _1992_/A _1984_/A VDD VSS sg13g2_nor2b_1
XFILLER_9_42 VDD VSS sg13g2_decap_8
X_1873_ _1872_/Y VDD _1884_/A VSS _1954_/S _1870_/B sg13g2_o21ai_1
XFILLER_30_763 VDD VSS sg13g2_decap_8
XFILLER_31_1043 VDD VSS sg13g2_decap_8
XFILLER_43_0 VDD VSS sg13g2_decap_8
XFILLER_9_1022 VDD VSS sg13g2_decap_8
XFILLER_85_936 VDD VSS sg13g2_decap_8
XFILLER_97_785 VDD VSS sg13g2_decap_8
XFILLER_97_796 VDD VSS sg13g2_fill_2
XFILLER_85_914 VDD VSS sg13g2_decap_8
XFILLER_96_273 VDD VSS sg13g2_decap_8
XFILLER_69_487 VDD VSS sg13g2_decap_8
X_2356_ _2356_/RESET_B VSS VDD _2356_/D _2356_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_111_595 VDD VSS sg13g2_decap_8
X_1307_ VDD _2183_/D _1307_/A VSS sg13g2_inv_1
XFILLER_84_435 VDD VSS sg13g2_decap_4
X_2295__129 VDD VSS _2295_/RESET_B sg13g2_tiehi
XFILLER_29_329 VDD VSS sg13g2_decap_8
X_2287_ _2287_/RESET_B VSS VDD _2287_/D _2287_/Q _2289_/CLK sg13g2_dfrbpq_1
X_1238_ _2092_/A _2093_/A _1238_/B VDD VSS sg13g2_nand2_1
XFILLER_38_863 VDD VSS sg13g2_decap_8
XFILLER_56_159 VDD VSS sg13g2_decap_8
XFILLER_71_118 VDD VSS sg13g2_decap_8
XFILLER_71_129 VDD VSS sg13g2_fill_1
XFILLER_65_682 VDD VSS sg13g2_decap_8
XFILLER_80_630 VDD VSS sg13g2_decap_8
X_2336__159 VDD VSS _2336_/RESET_B sg13g2_tiehi
XFILLER_53_866 VDD VSS sg13g2_decap_8
XFILLER_25_546 VDD VSS sg13g2_decap_8
XFILLER_44_28 VDD VSS sg13g2_decap_8
XFILLER_80_685 VDD VSS sg13g2_decap_8
XFILLER_80_696 VDD VSS sg13g2_fill_2
XFILLER_40_505 VDD VSS sg13g2_decap_8
XFILLER_100_56 VDD VSS sg13g2_decap_8
XFILLER_21_763 VDD VSS sg13g2_decap_8
XFILLER_20_273 VDD VSS sg13g2_decap_8
XFILLER_109_21 VDD VSS sg13g2_decap_8
XFILLER_4_406 VDD VSS sg13g2_decap_8
XFILLER_107_835 VDD VSS sg13g2_decap_8
XFILLER_106_312 VDD VSS sg13g2_decap_8
XFILLER_69_14 VDD VSS sg13g2_decap_8
XFILLER_109_98 VDD VSS sg13g2_decap_8
XFILLER_0_623 VDD VSS sg13g2_decap_8
XFILLER_88_774 VDD VSS sg13g2_decap_8
XFILLER_76_914 VDD VSS sg13g2_decap_4
XFILLER_87_262 VDD VSS sg13g2_decap_8
XFILLER_85_35 VDD VSS sg13g2_decap_8
XFILLER_102_595 VDD VSS sg13g2_decap_8
XFILLER_48_638 VDD VSS sg13g2_decap_8
XFILLER_75_479 VDD VSS sg13g2_decap_8
XFILLER_47_148 VDD VSS sg13g2_fill_1
XFILLER_84_980 VDD VSS sg13g2_decap_8
XFILLER_56_693 VDD VSS sg13g2_decap_8
XFILLER_44_811 VDD VSS sg13g2_decap_8
XFILLER_29_896 VDD VSS sg13g2_decap_8
XFILLER_18_84 VDD VSS sg13g2_decap_8
XFILLER_16_546 VDD VSS sg13g2_decap_8
XFILLER_43_343 VDD VSS sg13g2_decap_8
XFILLER_70_140 VDD VSS sg13g2_decap_8
XFILLER_54_1043 VDD VSS sg13g2_decap_8
XFILLER_12_763 VDD VSS sg13g2_decap_8
XFILLER_11_273 VDD VSS sg13g2_decap_8
XFILLER_8_756 VDD VSS sg13g2_decap_8
XFILLER_7_266 VDD VSS sg13g2_decap_8
XFILLER_109_161 VDD VSS sg13g2_decap_8
XFILLER_112_315 VDD VSS sg13g2_decap_8
XFILLER_4_973 VDD VSS sg13g2_decap_8
X_2210_ _2210_/RESET_B VSS VDD _2210_/D _2210_/Q clkload4/A sg13g2_dfrbpq_1
XFILLER_3_483 VDD VSS sg13g2_decap_8
XFILLER_79_785 VDD VSS sg13g2_decap_8
XFILLER_61_1047 VDD VSS sg13g2_decap_8
XFILLER_67_903 VDD VSS sg13g2_decap_8
XFILLER_39_605 VDD VSS sg13g2_decap_8
X_2141_ VDD VSS _2124_/B _2120_/A _2140_/X hold375/X _2143_/A _2124_/Y sg13g2_a221oi_1
XFILLER_78_295 VDD VSS sg13g2_decap_8
XFILLER_66_413 VDD VSS sg13g2_decap_4
XFILLER_66_435 VDD VSS sg13g2_decap_8
XFILLER_38_126 VDD VSS sg13g2_decap_8
XFILLER_82_928 VDD VSS sg13g2_decap_8
XFILLER_94_788 VDD VSS sg13g2_fill_1
X_2072_ _2339_/D _2072_/A _2072_/B VDD VSS sg13g2_nand2_1
XFILLER_81_405 VDD VSS sg13g2_decap_8
XFILLER_35_833 VDD VSS sg13g2_decap_8
XFILLER_53_118 VDD VSS sg13g2_decap_4
XFILLER_90_961 VDD VSS sg13g2_fill_2
XFILLER_34_343 VDD VSS sg13g2_decap_8
XFILLER_46_192 VDD VSS sg13g2_decap_8
XFILLER_90_994 VDD VSS sg13g2_decap_8
X_2216__108 VDD VSS _2216_/RESET_B sg13g2_tiehi
X_2190__160 VDD VSS _2190_/RESET_B sg13g2_tiehi
X_1925_ _1985_/A _1985_/B _1978_/A VDD VSS sg13g2_nor2_1
XFILLER_30_560 VDD VSS sg13g2_decap_8
X_1856_ _1952_/A _1856_/A _1856_/B VDD VSS sg13g2_xnor2_1
X_1787_ _1912_/B _2214_/Q _2222_/Q VDD VSS sg13g2_xnor2_1
Xfanout5 _2037_/A _2074_/A VDD VSS sg13g2_buf_1
XFILLER_104_827 VDD VSS sg13g2_decap_8
XFILLER_103_348 VDD VSS sg13g2_decap_8
XFILLER_39_28 VDD VSS sg13g2_decap_8
XFILLER_112_882 VDD VSS sg13g2_decap_8
X_2339_ _2339_/RESET_B VSS VDD _2339_/D _2339_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_84_221 VDD VSS sg13g2_fill_1
XFILLER_69_295 VDD VSS sg13g2_decap_8
XFILLER_58_936 VDD VSS sg13g2_decap_8
XFILLER_29_126 VDD VSS sg13g2_decap_8
XFILLER_85_777 VDD VSS sg13g2_decap_8
XFILLER_111_392 VDD VSS sg13g2_decap_8
XFILLER_57_446 VDD VSS sg13g2_decap_8
XFILLER_38_660 VDD VSS sg13g2_decap_8
XFILLER_26_833 VDD VSS sg13g2_decap_8
XFILLER_55_49 VDD VSS sg13g2_decap_8
XFILLER_77_1021 VDD VSS sg13g2_decap_8
XFILLER_25_343 VDD VSS sg13g2_decap_8
XFILLER_80_460 VDD VSS sg13g2_decap_8
XFILLER_38_1038 VDD VSS sg13g2_decap_8
XFILLER_41_825 VDD VSS sg13g2_decap_8
XFILLER_111_77 VDD VSS sg13g2_decap_8
XFILLER_40_335 VDD VSS sg13g2_decap_8
XFILLER_52_195 VDD VSS sg13g2_decap_8
XFILLER_21_560 VDD VSS sg13g2_decap_8
XFILLER_101_1041 VDD VSS sg13g2_decap_8
XFILLER_107_632 VDD VSS sg13g2_decap_8
XFILLER_4_203 VDD VSS sg13g2_decap_8
XFILLER_106_175 VDD VSS sg13g2_decap_8
XFILLER_20_63 VDD VSS sg13g2_decap_8
XFILLER_1_910 VDD VSS sg13g2_decap_8
XFILLER_84_1058 VDD VSS sg13g2_fill_2
XFILLER_0_420 VDD VSS sg13g2_decap_8
XFILLER_96_56 VDD VSS sg13g2_decap_8
XFILLER_1_987 VDD VSS sg13g2_decap_8
XFILLER_48_402 VDD VSS sg13g2_decap_8
XFILLER_88_582 VDD VSS sg13g2_decap_8
XFILLER_0_497 VDD VSS sg13g2_decap_8
XFILLER_76_755 VDD VSS sg13g2_decap_8
XFILLER_75_243 VDD VSS sg13g2_decap_8
XFILLER_90_202 VDD VSS sg13g2_decap_8
XFILLER_90_213 VDD VSS sg13g2_fill_1
XFILLER_90_235 VDD VSS sg13g2_decap_8
XFILLER_29_693 VDD VSS sg13g2_decap_8
XFILLER_56_490 VDD VSS sg13g2_decap_8
XFILLER_17_833 VDD VSS sg13g2_decap_8
XFILLER_91_1007 VDD VSS sg13g2_decap_8
XFILLER_72_983 VDD VSS sg13g2_decap_8
XFILLER_71_460 VDD VSS sg13g2_decap_8
XFILLER_16_343 VDD VSS sg13g2_decap_8
XFILLER_43_140 VDD VSS sg13g2_decap_8
XFILLER_32_847 VDD VSS sg13g2_decap_8
XFILLER_31_357 VDD VSS sg13g2_decap_8
XFILLER_84_7 VDD VSS sg13g2_decap_8
XFILLER_12_560 VDD VSS sg13g2_decap_8
XFILLER_61_70 VDD VSS sg13g2_decap_8
X_1710_ _1710_/Y _1720_/A _1710_/B VDD VSS sg13g2_nand2_1
XFILLER_8_553 VDD VSS sg13g2_decap_8
XFILLER_61_81 VDD VSS sg13g2_fill_1
X_1641_ _1688_/B _1641_/B _2307_/D VDD VSS sg13g2_and2_1
XFILLER_6_21 VDD VSS sg13g2_decap_8
XFILLER_99_836 VDD VSS sg13g2_decap_8
X_1572_ VSS VDD _1573_/A1 _1829_/A _1572_/Y _1523_/B sg13g2_a21oi_1
XFILLER_6_98 VDD VSS sg13g2_decap_8
XFILLER_4_770 VDD VSS sg13g2_decap_8
XFILLER_98_346 VDD VSS sg13g2_decap_8
XFILLER_112_112 VDD VSS sg13g2_decap_8
XFILLER_3_280 VDD VSS sg13g2_decap_8
XFILLER_100_307 VDD VSS sg13g2_decap_8
XFILLER_112_189 VDD VSS sg13g2_decap_8
XFILLER_6_1036 VDD VSS sg13g2_decap_8
X_2124_ _2124_/A _2124_/B _2124_/Y VDD VSS sg13g2_nor2_1
XFILLER_94_563 VDD VSS sg13g2_decap_4
XFILLER_39_457 VDD VSS sg13g2_decap_8
XFILLER_67_788 VDD VSS sg13g2_decap_4
XFILLER_66_287 VDD VSS sg13g2_decap_8
XFILLER_82_758 VDD VSS sg13g2_decap_8
X_2055_ _2055_/Y _2079_/S _2055_/B VDD VSS sg13g2_nand2_1
XFILLER_35_630 VDD VSS sg13g2_decap_8
XFILLER_34_140 VDD VSS sg13g2_decap_8
XFILLER_90_780 VDD VSS sg13g2_decap_8
XFILLER_50_611 VDD VSS sg13g2_decap_8
XFILLER_23_847 VDD VSS sg13g2_decap_8
XFILLER_22_357 VDD VSS sg13g2_decap_8
X_1908_ VDD _1908_/Y _1908_/A VSS sg13g2_inv_1
XFILLER_108_429 VDD VSS sg13g2_decap_8
X_1839_ _2245_/Q _2204_/Q _1839_/Y VDD VSS sg13g2_nor2b_1
Xhold520 _2275_/Q VDD VSS hold520/X sg13g2_dlygate4sd3_1
Xhold531 _1513_/Y VDD VSS _2271_/D sg13g2_dlygate4sd3_1
XFILLER_2_707 VDD VSS sg13g2_decap_8
Xhold542 _2296_/Q VDD VSS hold542/X sg13g2_dlygate4sd3_1
Xhold553 _1621_/Y VDD VSS _2293_/D sg13g2_dlygate4sd3_1
XFILLER_89_335 VDD VSS sg13g2_decap_8
XFILLER_103_112 VDD VSS sg13g2_decap_8
Xhold564 _2373_/Q VDD VSS hold564/X sg13g2_dlygate4sd3_1
XFILLER_1_217 VDD VSS sg13g2_decap_8
XFILLER_104_668 VDD VSS sg13g2_decap_8
XFILLER_58_700 VDD VSS sg13g2_decap_8
XFILLER_98_891 VDD VSS sg13g2_decap_8
XFILLER_103_189 VDD VSS sg13g2_decap_8
XFILLER_106_77 VDD VSS sg13g2_decap_8
XFILLER_73_714 VDD VSS sg13g2_decap_8
XFILLER_58_788 VDD VSS sg13g2_decap_8
XFILLER_57_276 VDD VSS sg13g2_decap_8
XFILLER_72_235 VDD VSS sg13g2_decap_4
XFILLER_82_14 VDD VSS sg13g2_decap_8
XFILLER_26_630 VDD VSS sg13g2_decap_8
XFILLER_54_983 VDD VSS sg13g2_decap_8
XFILLER_60_419 VDD VSS sg13g2_fill_2
XFILLER_25_140 VDD VSS sg13g2_decap_8
XFILLER_41_622 VDD VSS sg13g2_decap_8
XFILLER_14_847 VDD VSS sg13g2_decap_8
XFILLER_80_290 VDD VSS sg13g2_decap_8
XFILLER_13_357 VDD VSS sg13g2_decap_8
XFILLER_15_63 VDD VSS sg13g2_decap_8
XFILLER_51_1024 VDD VSS sg13g2_decap_8
XFILLER_41_699 VDD VSS sg13g2_decap_8
XFILLER_40_154 VDD VSS sg13g2_decap_8
X_2169__202 VDD VSS _2169_/RESET_B sg13g2_tiehi
XFILLER_12_1008 VDD VSS sg13g2_decap_8
XFILLER_108_941 VDD VSS sg13g2_decap_8
XFILLER_110_0 VDD VSS sg13g2_decap_8
XFILLER_31_84 VDD VSS sg13g2_decap_8
XFILLER_107_451 VDD VSS sg13g2_decap_8
XFILLER_5_567 VDD VSS sg13g2_decap_8
XFILLER_68_519 VDD VSS sg13g2_fill_2
XFILLER_68_508 VDD VSS sg13g2_decap_8
XFILLER_110_627 VDD VSS sg13g2_decap_8
XFILLER_89_880 VDD VSS sg13g2_decap_8
XFILLER_49_711 VDD VSS sg13g2_decap_8
XFILLER_1_784 VDD VSS sg13g2_decap_8
XFILLER_95_349 VDD VSS sg13g2_decap_4
XFILLER_37_917 VDD VSS sg13g2_decap_8
XFILLER_49_755 VDD VSS sg13g2_decap_8
XFILLER_0_294 VDD VSS sg13g2_decap_8
XFILLER_76_596 VDD VSS sg13g2_decap_8
XFILLER_64_725 VDD VSS sg13g2_decap_8
XFILLER_36_427 VDD VSS sg13g2_decap_8
XFILLER_17_630 VDD VSS sg13g2_decap_8
XFILLER_29_490 VDD VSS sg13g2_decap_8
XFILLER_91_577 VDD VSS sg13g2_decap_8
XFILLER_45_961 VDD VSS sg13g2_decap_8
XFILLER_16_140 VDD VSS sg13g2_decap_8
XFILLER_72_780 VDD VSS sg13g2_decap_8
XFILLER_60_942 VDD VSS sg13g2_decap_8
XFILLER_44_460 VDD VSS sg13g2_decap_8
XFILLER_108_1025 VDD VSS sg13g2_decap_8
XFILLER_32_644 VDD VSS sg13g2_decap_8
XFILLER_31_154 VDD VSS sg13g2_decap_8
XFILLER_9_840 VDD VSS sg13g2_decap_8
XFILLER_8_350 VDD VSS sg13g2_decap_8
X_1624_ _1624_/Y _1634_/A _1624_/B VDD VSS sg13g2_nand2_1
XFILLER_67_1053 VDD VSS sg13g2_decap_8
XFILLER_28_1015 VDD VSS sg13g2_decap_8
X_1555_ _1576_/A _1555_/B _2278_/D VDD VSS sg13g2_nor2_1
XFILLER_99_666 VDD VSS sg13g2_decap_8
X_1486_ VSS VDD _2093_/B hold392/X _1486_/Y _2101_/A sg13g2_a21oi_1
XFILLER_39_210 VDD VSS sg13g2_decap_8
XFILLER_86_349 VDD VSS sg13g2_decap_8
XFILLER_100_126 VDD VSS sg13g2_decap_8
XFILLER_28_917 VDD VSS sg13g2_decap_8
XFILLER_67_574 VDD VSS sg13g2_decap_8
XFILLER_55_769 VDD VSS sg13g2_decap_8
XFILLER_54_235 VDD VSS sg13g2_fill_1
Xclkbuf_leaf_19_clk clkbuf_leaf_0_clk/A clkload3/A VDD VSS sg13g2_buf_8
XFILLER_27_427 VDD VSS sg13g2_decap_8
X_2107_ _2107_/B1 VDD _2107_/Y VSS _1220_/A _2103_/Y sg13g2_o21ai_1
X_2038_ _2014_/X _2017_/B _2089_/S _2038_/X VDD VSS sg13g2_mux2_1
XFILLER_82_555 VDD VSS sg13g2_decap_8
XFILLER_70_717 VDD VSS sg13g2_decap_8
XFILLER_54_268 VDD VSS sg13g2_decap_8
XFILLER_42_419 VDD VSS sg13g2_decap_8
XFILLER_74_1024 VDD VSS sg13g2_decap_8
XFILLER_36_994 VDD VSS sg13g2_decap_8
XFILLER_51_975 VDD VSS sg13g2_decap_8
XFILLER_35_1008 VDD VSS sg13g2_decap_8
XFILLER_23_644 VDD VSS sg13g2_decap_8
XFILLER_50_430 VDD VSS sg13g2_decap_8
XFILLER_22_154 VDD VSS sg13g2_decap_8
XFILLER_109_749 VDD VSS sg13g2_decap_8
XFILLER_2_504 VDD VSS sg13g2_decap_8
Xhold361 _1290_/Y VDD VSS _1291_/A sg13g2_dlygate4sd3_1
XFILLER_104_421 VDD VSS sg13g2_fill_1
Xhold350 _2259_/Q VDD VSS _1194_/A sg13g2_dlygate4sd3_1
XFILLER_105_966 VDD VSS sg13g2_decap_8
XFILLER_78_806 VDD VSS sg13g2_decap_8
XFILLER_104_465 VDD VSS sg13g2_decap_8
XFILLER_89_154 VDD VSS sg13g2_decap_8
XFILLER_77_14 VDD VSS sg13g2_decap_8
Xhold394 _2164_/Q VDD VSS hold394/X sg13g2_dlygate4sd3_1
Xhold383 _2185_/Q VDD VSS hold383/X sg13g2_dlygate4sd3_1
Xhold372 _1225_/X VDD VSS _2359_/D sg13g2_dlygate4sd3_1
XFILLER_104_498 VDD VSS sg13g2_decap_8
XFILLER_92_319 VDD VSS sg13g2_decap_8
XFILLER_58_563 VDD VSS sg13g2_decap_8
XFILLER_46_703 VDD VSS sg13g2_decap_8
XFILLER_46_714 VDD VSS sg13g2_fill_1
XFILLER_19_917 VDD VSS sg13g2_decap_8
XFILLER_100_682 VDD VSS sg13g2_decap_8
XFILLER_93_35 VDD VSS sg13g2_decap_8
XFILLER_46_747 VDD VSS sg13g2_decap_8
XFILLER_18_427 VDD VSS sg13g2_decap_8
XFILLER_61_728 VDD VSS sg13g2_decap_8
XFILLER_42_931 VDD VSS sg13g2_decap_8
XFILLER_27_994 VDD VSS sg13g2_decap_8
XFILLER_26_84 VDD VSS sg13g2_decap_8
XFILLER_60_249 VDD VSS sg13g2_decap_8
XFILLER_14_644 VDD VSS sg13g2_decap_8
XFILLER_41_430 VDD VSS sg13g2_decap_8
XFILLER_13_154 VDD VSS sg13g2_decap_8
XFILLER_9_147 VDD VSS sg13g2_decap_8
XFILLER_10_861 VDD VSS sg13g2_decap_8
XFILLER_6_854 VDD VSS sg13g2_decap_8
XFILLER_5_364 VDD VSS sg13g2_decap_8
XFILLER_47_7 VDD VSS sg13g2_decap_8
XFILLER_111_903 VDD VSS sg13g2_decap_8
X_1340_ _1340_/Y _1342_/B1 hold366/X _1342_/A2 _2333_/Q VDD VSS sg13g2_a22oi_1
XFILLER_69_839 VDD VSS sg13g2_fill_1
XFILLER_110_424 VDD VSS sg13g2_decap_8
XFILLER_68_305 VDD VSS sg13g2_decap_8
X_1271_ VDD _2165_/D _1271_/A VSS sg13g2_inv_1
XFILLER_96_658 VDD VSS sg13g2_decap_8
XFILLER_3_77 VDD VSS sg13g2_decap_8
XFILLER_1_581 VDD VSS sg13g2_decap_8
XFILLER_49_530 VDD VSS sg13g2_decap_8
XFILLER_95_168 VDD VSS sg13g2_decap_8
XFILLER_37_714 VDD VSS sg13g2_decap_8
XFILLER_67_91 VDD VSS sg13g2_decap_8
XFILLER_64_522 VDD VSS sg13g2_decap_8
XFILLER_36_224 VDD VSS sg13g2_decap_8
XFILLER_97_1057 VDD VSS sg13g2_decap_4
XFILLER_91_341 VDD VSS sg13g2_decap_8
XFILLER_58_1019 VDD VSS sg13g2_fill_1
XFILLER_58_1008 VDD VSS sg13g2_decap_8
XFILLER_91_396 VDD VSS sg13g2_decap_8
XFILLER_33_931 VDD VSS sg13g2_decap_8
XFILLER_64_599 VDD VSS sg13g2_decap_8
XFILLER_18_994 VDD VSS sg13g2_decap_8
XFILLER_51_216 VDD VSS sg13g2_decap_8
XFILLER_32_441 VDD VSS sg13g2_decap_8
XFILLER_20_658 VDD VSS sg13g2_decap_8
XFILLER_73_0 VDD VSS sg13g2_decap_8
X_2310__290 VDD VSS _2310_/RESET_B sg13g2_tiehi
Xclkbuf_leaf_8_clk clkbuf_leaf_9_clk/A _2369_/CLK VDD VSS sg13g2_buf_8
X_1607_ _1612_/A _1607_/A _1618_/A VDD VSS sg13g2_xnor2_1
X_1538_ _1537_/Y VDD _1538_/Y VSS _1580_/A1 _2204_/Q sg13g2_o21ai_1
XFILLER_59_305 VDD VSS sg13g2_fill_2
XFILLER_80_1050 VDD VSS sg13g2_decap_8
XFILLER_87_658 VDD VSS sg13g2_decap_4
X_1469_ VSS VDD _1200_/Y _1481_/A2 _2253_/D _1468_/Y sg13g2_a21oi_1
XFILLER_47_28 VDD VSS sg13g2_decap_8
XFILLER_101_479 VDD VSS sg13g2_decap_8
XFILLER_86_157 VDD VSS sg13g2_decap_8
XFILLER_68_883 VDD VSS sg13g2_decap_8
XFILLER_28_714 VDD VSS sg13g2_decap_8
XFILLER_110_991 VDD VSS sg13g2_decap_8
XFILLER_41_1056 VDD VSS sg13g2_decap_4
XFILLER_55_522 VDD VSS sg13g2_decap_8
XFILLER_27_224 VDD VSS sg13g2_decap_8
XFILLER_83_864 VDD VSS sg13g2_decap_8
XFILLER_103_56 VDD VSS sg13g2_decap_8
XFILLER_24_931 VDD VSS sg13g2_decap_8
XFILLER_55_588 VDD VSS sg13g2_decap_8
XFILLER_36_791 VDD VSS sg13g2_decap_8
XFILLER_63_49 VDD VSS sg13g2_decap_8
XFILLER_42_205 VDD VSS sg13g2_decap_8
XFILLER_23_441 VDD VSS sg13g2_decap_8
XFILLER_42_238 VDD VSS sg13g2_decap_8
XFILLER_51_772 VDD VSS sg13g2_decap_8
XFILLER_11_658 VDD VSS sg13g2_decap_8
XFILLER_10_168 VDD VSS sg13g2_decap_8
XFILLER_109_546 VDD VSS sg13g2_decap_8
XFILLER_12_42 VDD VSS sg13g2_decap_8
XFILLER_88_35 VDD VSS sg13g2_decap_8
XFILLER_2_301 VDD VSS sg13g2_decap_8
XFILLER_105_763 VDD VSS sg13g2_decap_8
XFILLER_3_868 VDD VSS sg13g2_decap_8
XFILLER_78_614 VDD VSS sg13g2_decap_8
XFILLER_104_273 VDD VSS sg13g2_decap_8
XFILLER_2_378 VDD VSS sg13g2_decap_8
XFILLER_93_628 VDD VSS sg13g2_decap_8
XFILLER_77_168 VDD VSS sg13g2_decap_8
XFILLER_92_105 VDD VSS sg13g2_decap_8
XFILLER_59_883 VDD VSS sg13g2_fill_2
XFILLER_19_714 VDD VSS sg13g2_decap_8
XFILLER_74_842 VDD VSS sg13g2_decap_8
XFILLER_59_894 VDD VSS sg13g2_decap_8
XFILLER_18_224 VDD VSS sg13g2_decap_8
XFILLER_73_330 VDD VSS sg13g2_decap_8
XFILLER_46_544 VDD VSS sg13g2_decap_8
XFILLER_2_1050 VDD VSS sg13g2_decap_8
XFILLER_34_728 VDD VSS sg13g2_decap_8
XFILLER_27_791 VDD VSS sg13g2_decap_8
XFILLER_61_536 VDD VSS sg13g2_decap_8
XFILLER_15_931 VDD VSS sg13g2_decap_8
XFILLER_14_441 VDD VSS sg13g2_decap_8
XFILLER_33_238 VDD VSS sg13g2_decap_8
XFILLER_18_1036 VDD VSS sg13g2_decap_8
XFILLER_30_945 VDD VSS sg13g2_decap_8
XIO_FILL_IO_WEST_4_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
XFILLER_6_651 VDD VSS sg13g2_decap_8
XFILLER_5_161 VDD VSS sg13g2_decap_8
XFILLER_97_923 VDD VSS sg13g2_decap_8
XFILLER_111_700 VDD VSS sg13g2_decap_8
X_2372_ _2372_/RESET_B VSS VDD _2372_/D _2372_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_69_614 VDD VSS sg13g2_decap_8
XFILLER_64_1056 VDD VSS sg13g2_decap_4
XFILLER_97_967 VDD VSS sg13g2_fill_1
X_1323_ VDD _2191_/D _1323_/A VSS sg13g2_inv_1
XFILLER_110_210 VDD VSS sg13g2_decap_8
XFILLER_96_455 VDD VSS sg13g2_decap_8
XFILLER_25_1029 VDD VSS sg13g2_decap_8
XFILLER_68_124 VDD VSS sg13g2_fill_2
XFILLER_111_777 VDD VSS sg13g2_decap_8
XFILLER_84_606 VDD VSS sg13g2_decap_8
XFILLER_83_105 VDD VSS sg13g2_decap_8
X_1254_ _2271_/Q _1510_/A _1255_/B VDD VSS _1510_/B sg13g2_nand3b_1
XFILLER_56_319 VDD VSS sg13g2_decap_8
XFILLER_110_287 VDD VSS sg13g2_decap_8
XFILLER_65_820 VDD VSS sg13g2_decap_8
XFILLER_37_511 VDD VSS sg13g2_decap_8
XFILLER_92_661 VDD VSS sg13g2_decap_8
XFILLER_91_171 VDD VSS sg13g2_decap_8
XFILLER_37_588 VDD VSS sg13g2_decap_8
XFILLER_25_728 VDD VSS sg13g2_decap_8
XFILLER_64_374 VDD VSS sg13g2_decap_8
XFILLER_91_182 VDD VSS sg13g2_fill_1
XFILLER_52_569 VDD VSS sg13g2_decap_8
XFILLER_18_791 VDD VSS sg13g2_decap_8
XFILLER_24_238 VDD VSS sg13g2_decap_8
XFILLER_71_1005 VDD VSS sg13g2_decap_8
XFILLER_21_945 VDD VSS sg13g2_decap_8
XFILLER_60_580 VDD VSS sg13g2_decap_8
XFILLER_20_455 VDD VSS sg13g2_decap_8
XFILLER_0_805 VDD VSS sg13g2_decap_8
XFILLER_102_700 VDD VSS sg13g2_decap_8
XFILLER_102_744 VDD VSS sg13g2_decap_4
XFILLER_87_444 VDD VSS sg13g2_decap_8
XFILLER_58_49 VDD VSS sg13g2_fill_2
XFILLER_59_124 VDD VSS sg13g2_decap_8
XFILLER_102_766 VDD VSS sg13g2_decap_8
XFILLER_74_105 VDD VSS sg13g2_decap_8
XFILLER_101_276 VDD VSS sg13g2_decap_8
XFILLER_68_680 VDD VSS sg13g2_decap_8
XFILLER_28_511 VDD VSS sg13g2_decap_8
XFILLER_56_864 VDD VSS sg13g2_decap_8
XFILLER_71_812 VDD VSS sg13g2_decap_8
XFILLER_28_588 VDD VSS sg13g2_decap_8
XFILLER_55_385 VDD VSS sg13g2_decap_8
XFILLER_16_728 VDD VSS sg13g2_decap_8
XFILLER_43_569 VDD VSS sg13g2_decap_8
XFILLER_15_238 VDD VSS sg13g2_decap_8
XFILLER_90_14 VDD VSS sg13g2_decap_8
XFILLER_12_945 VDD VSS sg13g2_decap_8
XFILLER_11_455 VDD VSS sg13g2_decap_8
XFILLER_8_938 VDD VSS sg13g2_decap_8
XFILLER_23_63 VDD VSS sg13g2_decap_8
XFILLER_109_310 VDD VSS sg13g2_fill_2
XFILLER_7_448 VDD VSS sg13g2_decap_8
XFILLER_109_354 VDD VSS sg13g2_decap_8
XFILLER_99_56 VDD VSS sg13g2_decap_8
XFILLER_3_0 VDD VSS sg13g2_decap_8
XFILLER_79_934 VDD VSS sg13g2_decap_4
XFILLER_3_665 VDD VSS sg13g2_decap_8
XFILLER_2_175 VDD VSS sg13g2_decap_8
XFILLER_79_989 VDD VSS sg13g2_decap_4
XFILLER_93_414 VDD VSS sg13g2_decap_8
XFILLER_66_606 VDD VSS sg13g2_decap_4
XFILLER_94_948 VDD VSS sg13g2_decap_8
XFILLER_47_831 VDD VSS sg13g2_decap_8
XFILLER_19_511 VDD VSS sg13g2_decap_8
XFILLER_111_1043 VDD VSS sg13g2_decap_8
XFILLER_73_171 VDD VSS sg13g2_decap_8
XFILLER_0_56 VDD VSS sg13g2_decap_8
XFILLER_19_588 VDD VSS sg13g2_decap_8
XFILLER_34_525 VDD VSS sg13g2_decap_8
X_2177__186 VDD VSS _2177_/RESET_B sg13g2_tiehi
XFILLER_62_878 VDD VSS sg13g2_decap_8
XFILLER_9_21 VDD VSS sg13g2_decap_8
X_1941_ VSS VDD _2048_/A _2003_/B _1992_/B _1939_/Y sg13g2_a21oi_1
XFILLER_30_742 VDD VSS sg13g2_decap_8
X_1872_ _1872_/Y _1954_/S _2086_/A VDD VSS sg13g2_nand2_1
XFILLER_70_1060 VDD VSS sg13g2_fill_1
XFILLER_80_91 VDD VSS sg13g2_decap_8
XFILLER_31_1022 VDD VSS sg13g2_decap_8
XFILLER_9_98 VDD VSS sg13g2_decap_8
XFILLER_69_400 VDD VSS sg13g2_decap_8
XFILLER_9_1001 VDD VSS sg13g2_decap_8
XFILLER_69_422 VDD VSS sg13g2_decap_8
X_2355_ _2355_/RESET_B VSS VDD _2355_/D _2355_/Q clkload2/A sg13g2_dfrbpq_1
XFILLER_36_0 VDD VSS sg13g2_decap_8
XFILLER_111_574 VDD VSS sg13g2_decap_8
X_1306_ _1306_/Y _1322_/B1 hold387/X _1322_/A2 _2347_/Q VDD VSS sg13g2_a22oi_1
XFILLER_97_764 VDD VSS sg13g2_decap_8
XFILLER_96_252 VDD VSS sg13g2_decap_8
XFILLER_84_403 VDD VSS sg13g2_fill_1
XFILLER_69_466 VDD VSS sg13g2_decap_8
XFILLER_29_308 VDD VSS sg13g2_decap_8
XFILLER_57_639 VDD VSS sg13g2_decap_8
XFILLER_56_138 VDD VSS sg13g2_decap_8
X_2286_ _2286_/RESET_B VSS VDD _2286_/D _2286_/Q _2289_/CLK sg13g2_dfrbpq_1
XFILLER_38_842 VDD VSS sg13g2_decap_8
X_1237_ _1236_/Y VDD _1237_/Y VSS _1235_/A _1409_/C sg13g2_o21ai_1
XFILLER_25_525 VDD VSS sg13g2_decap_8
XFILLER_37_385 VDD VSS sg13g2_decap_8
XFILLER_52_300 VDD VSS sg13g2_decap_8
XFILLER_92_491 VDD VSS sg13g2_decap_8
XFILLER_53_845 VDD VSS sg13g2_decap_8
XFILLER_64_171 VDD VSS sg13g2_fill_1
XFILLER_80_664 VDD VSS sg13g2_decap_8
XFILLER_100_35 VDD VSS sg13g2_decap_8
XFILLER_21_742 VDD VSS sg13g2_decap_8
XIO_BOND_rst_n_pad rst_n_PAD bondpad_70x70
XFILLER_20_252 VDD VSS sg13g2_decap_8
XFILLER_107_814 VDD VSS sg13g2_decap_8
XFILLER_109_77 VDD VSS sg13g2_decap_8
XFILLER_106_379 VDD VSS sg13g2_decap_8
XFILLER_0_602 VDD VSS sg13g2_decap_8
XFILLER_85_14 VDD VSS sg13g2_decap_8
XFILLER_48_617 VDD VSS sg13g2_decap_8
XFILLER_0_679 VDD VSS sg13g2_decap_8
XFILLER_102_574 VDD VSS sg13g2_decap_8
XFILLER_75_425 VDD VSS sg13g2_decap_8
XFILLER_75_447 VDD VSS sg13g2_fill_2
XFILLER_75_458 VDD VSS sg13g2_decap_8
XFILLER_90_417 VDD VSS sg13g2_decap_8
XFILLER_56_683 VDD VSS sg13g2_decap_4
XFILLER_56_672 VDD VSS sg13g2_decap_8
XFILLER_29_875 VDD VSS sg13g2_decap_8
XFILLER_16_525 VDD VSS sg13g2_decap_8
XFILLER_18_63 VDD VSS sg13g2_decap_8
XFILLER_83_480 VDD VSS sg13g2_decap_8
XFILLER_55_182 VDD VSS sg13g2_decap_8
XFILLER_28_385 VDD VSS sg13g2_decap_8
XFILLER_71_675 VDD VSS sg13g2_decap_8
XFILLER_54_1011 VDD VSS sg13g2_decap_4
XFILLER_31_539 VDD VSS sg13g2_decap_8
XFILLER_43_399 VDD VSS sg13g2_decap_8
XFILLER_12_742 VDD VSS sg13g2_decap_8
XFILLER_34_84 VDD VSS sg13g2_decap_8
XFILLER_11_252 VDD VSS sg13g2_decap_8
XFILLER_8_735 VDD VSS sg13g2_decap_8
XFILLER_109_140 VDD VSS sg13g2_decap_8
XFILLER_7_245 VDD VSS sg13g2_decap_8
XFILLER_50_72 VDD VSS sg13g2_decap_8
XFILLER_109_184 VDD VSS sg13g2_fill_1
XFILLER_4_952 VDD VSS sg13g2_decap_8
XFILLER_98_539 VDD VSS sg13g2_decap_8
XFILLER_3_462 VDD VSS sg13g2_decap_8
XFILLER_79_764 VDD VSS sg13g2_decap_8
XFILLER_61_1026 VDD VSS sg13g2_decap_8
XFILLER_94_734 VDD VSS sg13g2_decap_4
X_2140_ _1510_/A _2201_/Q _2193_/Q _2185_/Q _2177_/Q _1510_/B _2140_/X VDD VSS sg13g2_mux4_1
XFILLER_78_285 VDD VSS sg13g2_decap_4
XFILLER_67_937 VDD VSS sg13g2_decap_4
XFILLER_38_105 VDD VSS sg13g2_decap_8
XFILLER_82_907 VDD VSS sg13g2_decap_8
X_2071_ _2071_/B _2071_/C _2071_/A _2072_/B VDD VSS sg13g2_nand3_1
XFILLER_93_233 VDD VSS sg13g2_fill_2
XFILLER_75_970 VDD VSS sg13g2_decap_8
XFILLER_93_277 VDD VSS sg13g2_decap_4
XFILLER_75_91 VDD VSS sg13g2_decap_8
XFILLER_35_812 VDD VSS sg13g2_decap_8
XFILLER_62_631 VDD VSS sg13g2_decap_8
XFILLER_19_385 VDD VSS sg13g2_decap_8
XFILLER_34_322 VDD VSS sg13g2_decap_8
XFILLER_90_973 VDD VSS sg13g2_decap_8
XFILLER_62_686 VDD VSS sg13g2_decap_8
XFILLER_50_826 VDD VSS sg13g2_decap_8
XFILLER_35_889 VDD VSS sg13g2_decap_8
XFILLER_61_185 VDD VSS sg13g2_decap_8
XFILLER_22_539 VDD VSS sg13g2_decap_8
XFILLER_34_399 VDD VSS sg13g2_decap_8
X_1924_ _1924_/B _1924_/A _1985_/B VDD VSS sg13g2_xor2_1
X_1855_ _1869_/A VDD _1954_/S VSS _2251_/Q _1208_/Y sg13g2_o21ai_1
X_1786_ VSS VDD _1900_/A _1900_/B _1912_/A _1779_/Y sg13g2_a21oi_1
X_2266__221 VDD VSS _2266_/RESET_B sg13g2_tiehi
XFILLER_104_806 VDD VSS sg13g2_decap_8
Xfanout6 _2054_/S _2069_/S VDD VSS sg13g2_buf_1
XFILLER_103_327 VDD VSS sg13g2_decap_8
XFILLER_112_861 VDD VSS sg13g2_decap_8
XFILLER_58_915 VDD VSS sg13g2_decap_8
X_2338_ _2338_/RESET_B VSS VDD _2338_/D _2338_/Q _2372_/CLK sg13g2_dfrbpq_1
XFILLER_111_371 VDD VSS sg13g2_decap_8
XFILLER_69_274 VDD VSS sg13g2_decap_8
XFILLER_58_959 VDD VSS sg13g2_fill_1
XFILLER_57_425 VDD VSS sg13g2_decap_8
XFILLER_29_105 VDD VSS sg13g2_decap_8
XFILLER_85_756 VDD VSS sg13g2_decap_8
XFILLER_84_255 VDD VSS sg13g2_fill_1
X_2269_ _2269_/RESET_B VSS VDD _2269_/D _2269_/Q _2365_/CLK sg13g2_dfrbpq_1
XFILLER_77_1000 VDD VSS sg13g2_decap_8
XFILLER_66_970 VDD VSS sg13g2_decap_8
XFILLER_26_812 VDD VSS sg13g2_decap_8
XFILLER_55_28 VDD VSS sg13g2_decap_8
XFILLER_84_299 VDD VSS sg13g2_decap_8
XFILLER_65_480 VDD VSS sg13g2_decap_8
XFILLER_25_322 VDD VSS sg13g2_decap_8
XFILLER_37_182 VDD VSS sg13g2_decap_8
XFILLER_111_56 VDD VSS sg13g2_decap_8
XFILLER_38_1017 VDD VSS sg13g2_decap_8
XFILLER_41_804 VDD VSS sg13g2_decap_8
XFILLER_26_889 VDD VSS sg13g2_decap_8
XFILLER_53_697 VDD VSS sg13g2_decap_8
XFILLER_13_539 VDD VSS sg13g2_decap_8
XFILLER_25_399 VDD VSS sg13g2_decap_8
XFILLER_40_314 VDD VSS sg13g2_decap_8
XFILLER_71_49 VDD VSS sg13g2_decap_8
XFILLER_14_1050 VDD VSS sg13g2_decap_8
XFILLER_107_611 VDD VSS sg13g2_decap_8
XFILLER_20_42 VDD VSS sg13g2_decap_8
XFILLER_5_749 VDD VSS sg13g2_decap_8
XFILLER_84_1037 VDD VSS sg13g2_decap_8
XFILLER_107_688 VDD VSS sg13g2_decap_8
XFILLER_106_154 VDD VSS sg13g2_decap_8
XFILLER_4_259 VDD VSS sg13g2_decap_8
XFILLER_96_35 VDD VSS sg13g2_decap_8
XFILLER_110_809 VDD VSS sg13g2_decap_8
XFILLER_88_561 VDD VSS sg13g2_decap_8
XFILLER_49_904 VDD VSS sg13g2_decap_8
XFILLER_1_966 VDD VSS sg13g2_decap_8
XFILLER_76_734 VDD VSS sg13g2_decap_8
XFILLER_102_382 VDD VSS sg13g2_decap_8
XFILLER_0_476 VDD VSS sg13g2_decap_8
XFILLER_75_222 VDD VSS sg13g2_decap_8
XFILLER_36_609 VDD VSS sg13g2_decap_8
XFILLER_29_84 VDD VSS sg13g2_decap_8
XFILLER_48_458 VDD VSS sg13g2_decap_4
XFILLER_64_929 VDD VSS sg13g2_decap_4
XFILLER_21_1043 VDD VSS sg13g2_decap_8
XFILLER_29_672 VDD VSS sg13g2_decap_8
XFILLER_17_812 VDD VSS sg13g2_decap_8
XFILLER_35_119 VDD VSS sg13g2_decap_8
XFILLER_91_759 VDD VSS sg13g2_decap_8
XFILLER_75_299 VDD VSS sg13g2_decap_8
XFILLER_44_620 VDD VSS sg13g2_decap_8
XFILLER_16_322 VDD VSS sg13g2_decap_8
XFILLER_28_182 VDD VSS sg13g2_decap_8
XFILLER_72_962 VDD VSS sg13g2_decap_8
XFILLER_17_889 VDD VSS sg13g2_decap_8
XFILLER_44_697 VDD VSS sg13g2_decap_8
XFILLER_32_826 VDD VSS sg13g2_decap_8
XFILLER_16_399 VDD VSS sg13g2_decap_8
XFILLER_31_336 VDD VSS sg13g2_decap_8
XFILLER_43_196 VDD VSS sg13g2_decap_8
XFILLER_77_7 VDD VSS sg13g2_decap_8
XFILLER_8_532 VDD VSS sg13g2_decap_8
X_1640_ _1674_/A hold518/X _1641_/B VDD VSS sg13g2_nor2b_1
X_1571_ VDD _1571_/Y _1571_/A VSS sg13g2_inv_1
XFILLER_99_815 VDD VSS sg13g2_decap_8
XFILLER_6_77 VDD VSS sg13g2_decap_8
XFILLER_98_325 VDD VSS sg13g2_decap_8
XFILLER_79_561 VDD VSS sg13g2_decap_8
XFILLER_112_168 VDD VSS sg13g2_decap_8
XFILLER_67_712 VDD VSS sg13g2_fill_1
XFILLER_6_1015 VDD VSS sg13g2_decap_8
XFILLER_94_542 VDD VSS sg13g2_decap_8
X_2123_ _2124_/A _2197_/Q _2189_/Q _2181_/Q _2173_/Q _2144_/S1 _2123_/X VDD VSS sg13g2_mux4_1
XFILLER_27_609 VDD VSS sg13g2_decap_8
XFILLER_39_436 VDD VSS sg13g2_decap_8
XFILLER_82_737 VDD VSS sg13g2_decap_8
XFILLER_81_203 VDD VSS sg13g2_decap_8
XFILLER_55_929 VDD VSS sg13g2_decap_8
XFILLER_48_981 VDD VSS sg13g2_decap_8
XFILLER_26_119 VDD VSS sg13g2_decap_8
X_2054_ _2048_/A _1936_/Y _2054_/S _2055_/B VDD VSS sg13g2_mux2_1
XFILLER_54_439 VDD VSS sg13g2_decap_8
XFILLER_19_182 VDD VSS sg13g2_decap_8
XFILLER_63_973 VDD VSS sg13g2_decap_8
XFILLER_35_686 VDD VSS sg13g2_decap_8
XFILLER_23_826 VDD VSS sg13g2_decap_8
XFILLER_37_1050 VDD VSS sg13g2_decap_8
XFILLER_22_336 VDD VSS sg13g2_decap_8
XFILLER_34_196 VDD VSS sg13g2_decap_8
XFILLER_50_678 VDD VSS sg13g2_decap_8
XFILLER_108_408 VDD VSS sg13g2_decap_8
X_1907_ _1907_/B _1907_/A _1908_/A VDD VSS sg13g2_xor2_1
X_1838_ _1905_/A _1921_/A _1860_/A VDD VSS sg13g2_nor2b_1
Xhold510 _1497_/Y VDD VSS _2267_/D sg13g2_dlygate4sd3_1
X_1769_ _1770_/B _1948_/A _1769_/B VDD VSS sg13g2_nand2_1
Xhold521 _2217_/Q VDD VSS _1386_/A sg13g2_dlygate4sd3_1
Xhold554 _2220_/Q VDD VSS hold554/X sg13g2_dlygate4sd3_1
Xhold543 _1635_/Y VDD VSS _1636_/B sg13g2_dlygate4sd3_1
Xhold532 _2295_/Q VDD VSS hold532/X sg13g2_dlygate4sd3_1
XFILLER_104_647 VDD VSS sg13g2_decap_8
Xhold565 _2372_/Q VDD VSS hold565/X sg13g2_dlygate4sd3_1
XFILLER_89_314 VDD VSS sg13g2_decap_8
XFILLER_98_870 VDD VSS sg13g2_decap_8
XFILLER_77_509 VDD VSS sg13g2_decap_8
XFILLER_103_168 VDD VSS sg13g2_decap_8
XFILLER_106_56 VDD VSS sg13g2_decap_8
XFILLER_44_1054 VDD VSS sg13g2_decap_8
XFILLER_57_200 VDD VSS sg13g2_decap_8
XFILLER_46_918 VDD VSS sg13g2_decap_8
XFILLER_57_222 VDD VSS sg13g2_fill_2
XFILLER_18_609 VDD VSS sg13g2_decap_8
XFILLER_66_49 VDD VSS sg13g2_decap_8
XFILLER_100_875 VDD VSS sg13g2_fill_2
XFILLER_85_575 VDD VSS sg13g2_decap_8
XFILLER_72_214 VDD VSS sg13g2_decap_8
XFILLER_17_119 VDD VSS sg13g2_decap_8
XFILLER_45_428 VDD VSS sg13g2_fill_2
XFILLER_54_962 VDD VSS sg13g2_decap_8
XFILLER_41_601 VDD VSS sg13g2_decap_8
XFILLER_26_686 VDD VSS sg13g2_decap_8
XFILLER_14_826 VDD VSS sg13g2_decap_8
XFILLER_13_336 VDD VSS sg13g2_decap_8
XFILLER_15_42 VDD VSS sg13g2_decap_8
XFILLER_40_133 VDD VSS sg13g2_decap_8
XFILLER_25_196 VDD VSS sg13g2_decap_8
XFILLER_51_1003 VDD VSS sg13g2_decap_8
XFILLER_41_678 VDD VSS sg13g2_decap_8
XFILLER_9_329 VDD VSS sg13g2_decap_8
XFILLER_108_920 VDD VSS sg13g2_decap_8
XFILLER_107_430 VDD VSS sg13g2_decap_8
XFILLER_5_546 VDD VSS sg13g2_decap_8
XFILLER_31_63 VDD VSS sg13g2_decap_8
XFILLER_108_997 VDD VSS sg13g2_decap_8
XFILLER_103_0 VDD VSS sg13g2_decap_8
XFILLER_110_606 VDD VSS sg13g2_decap_8
XFILLER_96_829 VDD VSS sg13g2_decap_8
XFILLER_1_763 VDD VSS sg13g2_decap_8
XFILLER_95_328 VDD VSS sg13g2_decap_8
XFILLER_0_273 VDD VSS sg13g2_decap_8
XFILLER_88_380 VDD VSS sg13g2_decap_8
XFILLER_48_244 VDD VSS sg13g2_decap_4
XFILLER_76_564 VDD VSS sg13g2_decap_8
XFILLER_64_704 VDD VSS sg13g2_decap_8
XFILLER_36_406 VDD VSS sg13g2_decap_8
XFILLER_45_940 VDD VSS sg13g2_decap_8
XFILLER_56_71 VDD VSS sg13g2_fill_1
XFILLER_48_288 VDD VSS sg13g2_decap_8
XFILLER_91_556 VDD VSS sg13g2_decap_8
XFILLER_63_269 VDD VSS sg13g2_decap_8
XFILLER_108_1004 VDD VSS sg13g2_decap_8
XFILLER_60_921 VDD VSS sg13g2_decap_8
XFILLER_32_623 VDD VSS sg13g2_decap_8
XFILLER_17_686 VDD VSS sg13g2_decap_8
XFILLER_71_280 VDD VSS sg13g2_decap_8
XFILLER_71_291 VDD VSS sg13g2_fill_2
XFILLER_72_70 VDD VSS sg13g2_decap_8
XFILLER_16_196 VDD VSS sg13g2_decap_8
XFILLER_31_133 VDD VSS sg13g2_decap_8
XFILLER_9_896 VDD VSS sg13g2_decap_8
XFILLER_67_1032 VDD VSS sg13g2_decap_8
XFILLER_67_1010 VDD VSS sg13g2_fill_2
X_1623_ _1624_/B _1623_/A _1628_/A VDD VSS sg13g2_xnor2_1
X_1554_ _1555_/B _1527_/Y _1553_/Y hold478/X _1527_/B VDD VSS sg13g2_a22oi_1
XFILLER_87_829 VDD VSS sg13g2_decap_8
XFILLER_98_133 VDD VSS sg13g2_decap_8
XIO_FILL_IO_EAST_2_0 IOVDD IOVSS VDD VSS sg13g2_Filler200
X_1485_ _1485_/Y _1485_/A _1487_/B VDD VSS sg13g2_nand2_1
XFILLER_86_328 VDD VSS sg13g2_decap_8
XFILLER_86_306 VDD VSS sg13g2_fill_2
XFILLER_100_105 VDD VSS sg13g2_decap_8
.ends

